`timescale 1ns / 1ps

module ROM_W21(
    input [12:0] addr,
    output reg [15:0] weight
    );
    
always @(*)
    case(addr)
13'd0:weight<=16'b0000000000010110  ;
13'd1:weight<=16'b1111111111011100   ;
13'd2:weight<=16'b0000000001101011   ;
13'd3:weight<=16'b0000000000101111   ;
13'd4:weight<=16'b1111111111110110   ;
13'd5:weight<=16'b0000000010010011   ;
13'd6:weight<=16'b1111111110011111   ;
13'd7:weight<=16'b0000000000001010   ;
13'd8:weight<=16'b1111111111010010   ;
13'd9:weight<=16'b1111111110010110   ;
13'd10:weight<=16'b0000000001100110   ;
13'd11:weight<=16'b0000000000110100   ;
13'd12:weight<=16'b1111111011010110   ;
13'd13:weight<=16'b1111111110001011   ;
13'd14:weight<=16'b0000000011001110   ;
13'd15:weight<=16'b0000000001101000   ;
13'd16:weight<=16'b0000000001010010   ;
13'd17:weight<=16'b0000000000100000   ;
13'd18:weight<=16'b1111111011011010   ;
13'd19:weight<=16'b0000000010010100   ;
13'd20:weight<=16'b0000000001101111   ;
13'd21:weight<=16'b1111111110000110   ;
13'd22:weight<=16'b1111111110100100   ;
13'd23:weight<=16'b0000000010000001   ;
13'd24:weight<=16'b1111111101100011   ;
13'd25:weight<=16'b1111111100111000   ;
13'd26:weight<=16'b0000000000010011   ;
13'd27:weight<=16'b0000000100000001   ;
13'd28:weight<=16'b0000000100010010   ;
13'd29:weight<=16'b1111111101010111   ;
13'd30:weight<=16'b0000000000101010   ;
13'd31:weight<=16'b0000000000000100   ;
13'd32:weight<=16'b0000000000100100   ;
13'd33:weight<=16'b0000000001000110   ;
13'd34:weight<=16'b0000000110011011   ;
13'd35:weight<=16'b1111111111101110   ;
13'd36:weight<=16'b1111111101000110   ;
13'd37:weight<=16'b1111111110110010   ;
13'd38:weight<=16'b0000000100001100   ;
13'd39:weight<=16'b1111111000011000   ;
13'd40:weight<=16'b1111111111011100   ;
13'd41:weight<=16'b0000000100000010   ;
13'd42:weight<=16'b1111111101100101   ;
13'd43:weight<=16'b0000000000001001   ;
13'd44:weight<=16'b1111111101010110   ;
13'd45:weight<=16'b0000000001010100   ;
13'd46:weight<=16'b0000000001000111   ;
13'd47:weight<=16'b1111111101110011   ;
13'd48:weight<=16'b0000000000101101   ;
13'd49:weight<=16'b0000000001101011   ;
13'd50:weight<=16'b0000000000010110   ;
13'd51:weight<=16'b1111111111011100   ;
13'd52:weight<=16'b0000000001101011   ;
13'd53:weight<=16'b0000000000101111   ;
13'd54:weight<=16'b1111111111110110   ;
13'd55:weight<=16'b0000000010010011   ;
13'd56:weight<=16'b1111111110011111   ;
13'd57:weight<=16'b0000000000001010   ;
13'd58:weight<=16'b1111111111010010   ;
13'd59:weight<=16'b1111111110010110   ;
13'd60:weight<=16'b0000000000000010   ;
13'd61:weight<=16'b1111111111111110   ;
13'd62:weight<=16'b1111111110001011   ;
13'd63:weight<=16'b0000000011000110   ;
13'd64:weight<=16'b1111111111101001   ;
13'd65:weight<=16'b1111111111111111   ;
13'd66:weight<=16'b1111111111101110   ;
13'd67:weight<=16'b0000000000100101   ;
13'd68:weight<=16'b1111111101110011   ;
13'd69:weight<=16'b0000000001100000   ;
13'd70:weight<=16'b0000000001101111   ;
13'd71:weight<=16'b1111111110000110   ;
13'd72:weight<=16'b1111111110100100   ;
13'd73:weight<=16'b0000000010000001   ;
13'd74:weight<=16'b1111111101100011   ;
13'd75:weight<=16'b1111111100111000   ;
13'd76:weight<=16'b0000000000010011   ;
13'd77:weight<=16'b0000000100000001   ;
13'd78:weight<=16'b0000000100010010   ;
13'd79:weight<=16'b1111111101010111   ;
13'd80:weight<=16'b0000000100000101   ;
13'd81:weight<=16'b0000000000100110   ;
13'd82:weight<=16'b0000000000110100   ;
13'd83:weight<=16'b0000000001100000   ;
13'd84:weight<=16'b0000000001111100   ;
13'd85:weight<=16'b0000000000101110   ;
13'd86:weight<=16'b1111111011111000   ;
13'd87:weight<=16'b1111111110111110   ;
13'd88:weight<=16'b1111111110101000   ;
13'd89:weight<=16'b1111111110110101   ;
13'd90:weight<=16'b1111111111011100   ;
13'd91:weight<=16'b0000000100000010   ;
13'd92:weight<=16'b1111111101100101   ;
13'd93:weight<=16'b0000000000001001   ;
13'd94:weight<=16'b1111111101010110   ;
13'd95:weight<=16'b0000000001010100   ;
13'd96:weight<=16'b0000000001000111   ;
13'd97:weight<=16'b1111111101110011   ;
13'd98:weight<=16'b0000000000101101   ;
13'd99:weight<=16'b0000000001101011   ;
13'd100:weight<=16'b1111111111100110   ;
13'd101:weight<=16'b0000000000010110   ;
13'd102:weight<=16'b0000000000001010   ;
13'd103:weight<=16'b1111111111101010   ;
13'd104:weight<=16'b0000000001000011   ;
13'd105:weight<=16'b1111111101111111   ;
13'd106:weight<=16'b0000000001011010   ;
13'd107:weight<=16'b1111111110101101   ;
13'd108:weight<=16'b1111111101011011   ;
13'd109:weight<=16'b0000000100101010   ;
13'd110:weight<=16'b0000000000000010   ;
13'd111:weight<=16'b1111111111111110   ;
13'd112:weight<=16'b1111111110001011   ;
13'd113:weight<=16'b0000000011000110   ;
13'd114:weight<=16'b1111111111101001   ;
13'd115:weight<=16'b1111111111111111   ;
13'd116:weight<=16'b1111111111101110   ;
13'd117:weight<=16'b0000000000100101   ;
13'd118:weight<=16'b1111111101110011   ;
13'd119:weight<=16'b0000000001100000   ;
13'd120:weight<=16'b0000000000010011   ;
13'd121:weight<=16'b1111111111010100   ;
13'd122:weight<=16'b0000000010100010   ;
13'd123:weight<=16'b1111111110101111   ;
13'd124:weight<=16'b0000000000000101   ;
13'd125:weight<=16'b0000000000001001   ;
13'd126:weight<=16'b0000000000000110   ;
13'd127:weight<=16'b1111111111000010   ;
13'd128:weight<=16'b1111111111101011   ;
13'd129:weight<=16'b0000000000010101   ;
13'd130:weight<=16'b0000000100000101   ;
13'd131:weight<=16'b0000000000100110   ;
13'd132:weight<=16'b0000000000110100   ;
13'd133:weight<=16'b0000000001100000   ;
13'd134:weight<=16'b0000000001111100   ;
13'd135:weight<=16'b0000000000101110   ;
13'd136:weight<=16'b1111111011111000   ;
13'd137:weight<=16'b1111111110111110   ;
13'd138:weight<=16'b1111111110101000   ;
13'd139:weight<=16'b1111111110110101   ;
13'd140:weight<=16'b0000000001101100   ;
13'd141:weight<=16'b1111111110111011   ;
13'd142:weight<=16'b0000000010001011   ;
13'd143:weight<=16'b0000000000001111   ;
13'd144:weight<=16'b0000000001101110   ;
13'd145:weight<=16'b1111111101110111   ;
13'd146:weight<=16'b1111111110100100   ;
13'd147:weight<=16'b0000000000001001   ;
13'd148:weight<=16'b1111111101110110   ;
13'd149:weight<=16'b0000000010000010   ;
13'd150:weight<=16'b1111111111100110   ;
13'd151:weight<=16'b0000000000010110   ;
13'd152:weight<=16'b0000000000001010   ;
13'd153:weight<=16'b1111111111101010   ;
13'd154:weight<=16'b0000000001000011   ;
13'd155:weight<=16'b1111111101111111   ;
13'd156:weight<=16'b0000000001011010   ;
13'd157:weight<=16'b1111111110101101   ;
13'd158:weight<=16'b1111111101011011   ;
13'd159:weight<=16'b0000000100101010   ;
13'd160:weight<=16'b1111111111101111   ;
13'd161:weight<=16'b0000000010000100   ;
13'd162:weight<=16'b1111111110000010   ;
13'd163:weight<=16'b0000000000111101   ;
13'd164:weight<=16'b1111111111000010   ;
13'd165:weight<=16'b1111111110111100   ;
13'd166:weight<=16'b0000000010100111   ;
13'd167:weight<=16'b1111111110110001   ;
13'd168:weight<=16'b1111111111001011   ;
13'd169:weight<=16'b0000000000101111   ;
13'd170:weight<=16'b0000000000010011   ;
13'd171:weight<=16'b1111111111010100   ;
13'd172:weight<=16'b0000000010100010   ;
13'd173:weight<=16'b1111111110101111   ;
13'd174:weight<=16'b0000000000000101   ;
13'd175:weight<=16'b0000000000001001   ;
13'd176:weight<=16'b0000000000000110   ;
13'd177:weight<=16'b1111111111000010   ;
13'd178:weight<=16'b1111111111101011   ;
13'd179:weight<=16'b0000000000010101   ;
13'd180:weight<=16'b0000000010110010   ;
13'd181:weight<=16'b0000000000011101   ;
13'd182:weight<=16'b1111111111001011   ;
13'd183:weight<=16'b1111111111100101   ;
13'd184:weight<=16'b1111111101100000   ;
13'd185:weight<=16'b0000000001110000   ;
13'd186:weight<=16'b0000000000111111   ;
13'd187:weight<=16'b0000000010100110   ;
13'd188:weight<=16'b1111111110010111   ;
13'd189:weight<=16'b1111111110100001   ;
13'd190:weight<=16'b0000000001101100   ;
13'd191:weight<=16'b1111111110111011   ;
13'd192:weight<=16'b0000000010001011   ;
13'd193:weight<=16'b0000000000001111   ;
13'd194:weight<=16'b0000000001101110   ;
13'd195:weight<=16'b1111111101110111   ;
13'd196:weight<=16'b1111111110100100   ;
13'd197:weight<=16'b0000000000001001   ;
13'd198:weight<=16'b1111111101110110   ;
13'd199:weight<=16'b0000000010000010   ;
13'd200:weight<=16'b1111111111000100   ;
13'd201:weight<=16'b1111111110000110   ;
13'd202:weight<=16'b0000000010010001   ;
13'd203:weight<=16'b0000000000000100   ;
13'd204:weight<=16'b0000000000000110   ;
13'd205:weight<=16'b1111111110110111   ;
13'd206:weight<=16'b0000000000010111   ;
13'd207:weight<=16'b0000000000100001   ;
13'd208:weight<=16'b0000000000000111   ;
13'd209:weight<=16'b0000000010000111   ;
13'd210:weight<=16'b1111111111101111   ;
13'd211:weight<=16'b0000000010000100   ;
13'd212:weight<=16'b1111111110000010   ;
13'd213:weight<=16'b0000000000111101   ;
13'd214:weight<=16'b1111111111000010   ;
13'd215:weight<=16'b1111111110111100   ;
13'd216:weight<=16'b0000000010100111   ;
13'd217:weight<=16'b1111111110110001   ;
13'd218:weight<=16'b1111111111001011   ;
13'd219:weight<=16'b0000000000101111   ;
13'd220:weight<=16'b1111111110000111   ;
13'd221:weight<=16'b0000000011001010   ;
13'd222:weight<=16'b1111111111110001   ;
13'd223:weight<=16'b1111111111001011   ;
13'd224:weight<=16'b1111111110111110   ;
13'd225:weight<=16'b0000000001110010   ;
13'd226:weight<=16'b0000000001011000   ;
13'd227:weight<=16'b0000000010010111   ;
13'd228:weight<=16'b1111111110000000   ;
13'd229:weight<=16'b1111111111101111   ;
13'd230:weight<=16'b0000000010110010   ;
13'd231:weight<=16'b0000000000011101   ;
13'd232:weight<=16'b1111111111001011   ;
13'd233:weight<=16'b1111111111100101   ;
13'd234:weight<=16'b1111111101100000   ;
13'd235:weight<=16'b0000000001110000   ;
13'd236:weight<=16'b0000000000111111   ;
13'd237:weight<=16'b0000000010100110   ;
13'd238:weight<=16'b1111111110010111   ;
13'd239:weight<=16'b1111111110100001   ;
13'd240:weight<=16'b0000000001011001   ;
13'd241:weight<=16'b1111111111010101   ;
13'd242:weight<=16'b0000000001001101   ;
13'd243:weight<=16'b1111111101110000   ;
13'd244:weight<=16'b0000000000110001   ;
13'd245:weight<=16'b1111111111011110   ;
13'd246:weight<=16'b0000000010011010   ;
13'd247:weight<=16'b0000000000111100   ;
13'd248:weight<=16'b1111111111000010   ;
13'd249:weight<=16'b1111111110100001   ;
13'd250:weight<=16'b1111111111000100   ;
13'd251:weight<=16'b1111111110000110   ;
13'd252:weight<=16'b0000000010010001   ;
13'd253:weight<=16'b0000000000000100   ;
13'd254:weight<=16'b0000000000000110   ;
13'd255:weight<=16'b1111111110110111   ;
13'd256:weight<=16'b0000000000010111   ;
13'd257:weight<=16'b0000000000100001   ;
13'd258:weight<=16'b0000000000000111   ;
13'd259:weight<=16'b0000000010000111   ;
13'd260:weight<=16'b1111111111100100   ;
13'd261:weight<=16'b0000000010111001   ;
13'd262:weight<=16'b1111111110010000   ;
13'd263:weight<=16'b1111111111110101   ;
13'd264:weight<=16'b1111111110100010   ;
13'd265:weight<=16'b0000000001001011   ;
13'd266:weight<=16'b0000000000110111   ;
13'd267:weight<=16'b0000000001011000   ;
13'd268:weight<=16'b1111111110011111   ;
13'd269:weight<=16'b0000000000100000   ;
13'd270:weight<=16'b1111111110000111   ;
13'd271:weight<=16'b0000000011001010   ;
13'd272:weight<=16'b1111111111110001   ;
13'd273:weight<=16'b1111111111001011   ;
13'd274:weight<=16'b1111111110111110   ;
13'd275:weight<=16'b0000000001110010   ;
13'd276:weight<=16'b0000000001011000   ;
13'd277:weight<=16'b0000000010010111   ;
13'd278:weight<=16'b1111111110000000   ;
13'd279:weight<=16'b1111111111101111   ;
13'd280:weight<=16'b1111111111101101   ;
13'd281:weight<=16'b0000000001010000   ;
13'd282:weight<=16'b0000000000011111   ;
13'd283:weight<=16'b1111111101000000   ;
13'd284:weight<=16'b0000000000010010   ;
13'd285:weight<=16'b1111111111101101   ;
13'd286:weight<=16'b1111111110000101   ;
13'd287:weight<=16'b0000000001000000   ;
13'd288:weight<=16'b1111111111110010   ;
13'd289:weight<=16'b0000000011010101   ;
13'd290:weight<=16'b0000000001011001   ;
13'd291:weight<=16'b1111111111010101   ;
13'd292:weight<=16'b0000000001001101   ;
13'd293:weight<=16'b1111111101110000   ;
13'd294:weight<=16'b0000000000110001   ;
13'd295:weight<=16'b1111111111011110   ;
13'd296:weight<=16'b0000000010011010   ;
13'd297:weight<=16'b0000000000111100   ;
13'd298:weight<=16'b1111111111000010   ;
13'd299:weight<=16'b1111111110100001   ;
13'd300:weight<=16'b1111111110011011   ;
13'd301:weight<=16'b1111111111001101   ;
13'd302:weight<=16'b1111111110101001   ;
13'd303:weight<=16'b1111111110010010   ;
13'd304:weight<=16'b0000000010000111   ;
13'd305:weight<=16'b1111111101111100   ;
13'd306:weight<=16'b1111111111010100   ;
13'd307:weight<=16'b0000000001110101   ;
13'd308:weight<=16'b1111111111100000   ;
13'd309:weight<=16'b0000000101001101   ;
13'd310:weight<=16'b1111111111100100   ;
13'd311:weight<=16'b0000000010111001   ;
13'd312:weight<=16'b1111111110010000   ;
13'd313:weight<=16'b1111111111110101   ;
13'd314:weight<=16'b1111111110100010   ;
13'd315:weight<=16'b0000000001001011   ;
13'd316:weight<=16'b0000000000110111   ;
13'd317:weight<=16'b0000000001011000   ;
13'd318:weight<=16'b1111111110011111   ;
13'd319:weight<=16'b0000000000100000   ;
13'd320:weight<=16'b1111111110100001   ;
13'd321:weight<=16'b0000000001101000   ;
13'd322:weight<=16'b1111111110001010   ;
13'd323:weight<=16'b1111111110100111   ;
13'd324:weight<=16'b1111111111100010   ;
13'd325:weight<=16'b0000000001001011   ;
13'd326:weight<=16'b1111111110000100   ;
13'd327:weight<=16'b0000000100001001   ;
13'd328:weight<=16'b1111111110101001   ;
13'd329:weight<=16'b0000000010011101   ;
13'd330:weight<=16'b1111111111101101   ;
13'd331:weight<=16'b0000000001010000   ;
13'd332:weight<=16'b0000000000011111   ;
13'd333:weight<=16'b1111111101000000   ;
13'd334:weight<=16'b0000000000010010   ;
13'd335:weight<=16'b1111111111101101   ;
13'd336:weight<=16'b1111111110000101   ;
13'd337:weight<=16'b0000000001000000   ;
13'd338:weight<=16'b1111111111110010   ;
13'd339:weight<=16'b0000000011010101   ;
13'd340:weight<=16'b0000000011000010   ;
13'd341:weight<=16'b0000000000001011   ;
13'd342:weight<=16'b0000000000010110   ;
13'd343:weight<=16'b1111111110111110   ;
13'd344:weight<=16'b1111111111000101   ;
13'd345:weight<=16'b1111111111100001   ;
13'd346:weight<=16'b1111111111011010   ;
13'd347:weight<=16'b1111111111000101   ;
13'd348:weight<=16'b1111111111011011   ;
13'd349:weight<=16'b0000000001100000   ;
13'd350:weight<=16'b1111111110011011   ;
13'd351:weight<=16'b1111111111001101   ;
13'd352:weight<=16'b1111111110101001   ;
13'd353:weight<=16'b1111111110010010   ;
13'd354:weight<=16'b0000000010000111   ;
13'd355:weight<=16'b1111111101111100   ;
13'd356:weight<=16'b1111111111010100   ;
13'd357:weight<=16'b0000000001110101   ;
13'd358:weight<=16'b1111111111100000   ;
13'd359:weight<=16'b0000000101001101   ;
13'd360:weight<=16'b0000000000100000   ;
13'd361:weight<=16'b0000000000110011   ;
13'd362:weight<=16'b1111111111010011   ;
13'd363:weight<=16'b1111111111010010   ;
13'd364:weight<=16'b1111111110101011   ;
13'd365:weight<=16'b1111111110111111   ;
13'd366:weight<=16'b1111111111101001   ;
13'd367:weight<=16'b0000000010011111   ;
13'd368:weight<=16'b0000000001111001   ;
13'd369:weight<=16'b1111111110111111   ;
13'd370:weight<=16'b1111111110100001   ;
13'd371:weight<=16'b0000000001101000   ;
13'd372:weight<=16'b1111111110001010   ;
13'd373:weight<=16'b1111111110100111   ;
13'd374:weight<=16'b1111111111100010   ;
13'd375:weight<=16'b0000000001001011   ;
13'd376:weight<=16'b1111111110000100   ;
13'd377:weight<=16'b0000000100001001   ;
13'd378:weight<=16'b1111111110101001   ;
13'd379:weight<=16'b0000000010011101   ;
13'd380:weight<=16'b0000000000000010   ;
13'd381:weight<=16'b0000000000101110   ;
13'd382:weight<=16'b0000000000100100   ;
13'd383:weight<=16'b1111111101000011   ;
13'd384:weight<=16'b1111111111000100   ;
13'd385:weight<=16'b0000000001010011   ;
13'd386:weight<=16'b0000000011000101   ;
13'd387:weight<=16'b0000000011110010   ;
13'd388:weight<=16'b1111111110001010   ;
13'd389:weight<=16'b1111111101111011   ;
13'd390:weight<=16'b0000000011000010   ;
13'd391:weight<=16'b0000000000001011   ;
13'd392:weight<=16'b0000000000010110   ;
13'd393:weight<=16'b1111111110111110   ;
13'd394:weight<=16'b1111111111000101   ;
13'd395:weight<=16'b1111111111100001   ;
13'd396:weight<=16'b1111111111011010   ;
13'd397:weight<=16'b1111111111000101   ;
13'd398:weight<=16'b1111111111011011   ;
13'd399:weight<=16'b0000000001100000   ;
13'd400:weight<=16'b0000000010001100   ;
13'd401:weight<=16'b0000000001011111   ;
13'd402:weight<=16'b1111111111100101   ;
13'd403:weight<=16'b1111111111100100   ;
13'd404:weight<=16'b1111111111100001   ;
13'd405:weight<=16'b1111111110110111   ;
13'd406:weight<=16'b1111111110101110   ;
13'd407:weight<=16'b0000000000010010   ;
13'd408:weight<=16'b0000000001100010   ;
13'd409:weight<=16'b1111111110101011   ;
13'd410:weight<=16'b0000000000100000   ;
13'd411:weight<=16'b0000000000110011   ;
13'd412:weight<=16'b1111111111010011   ;
13'd413:weight<=16'b1111111111010010   ;
13'd414:weight<=16'b1111111110101011   ;
13'd415:weight<=16'b1111111110111111   ;
13'd416:weight<=16'b1111111111101001   ;
13'd417:weight<=16'b0000000010011111   ;
13'd418:weight<=16'b0000000001111001   ;
13'd419:weight<=16'b1111111110111111   ;
13'd420:weight<=16'b0000000010100010   ;
13'd421:weight<=16'b0000000001100001   ;
13'd422:weight<=16'b1111111101001011   ;
13'd423:weight<=16'b1111111111000010   ;
13'd424:weight<=16'b1111111101111111   ;
13'd425:weight<=16'b0000000001010000   ;
13'd426:weight<=16'b0000000000111010   ;
13'd427:weight<=16'b0000000100100000   ;
13'd428:weight<=16'b0000000000001000   ;
13'd429:weight<=16'b1111111101010010   ;
13'd430:weight<=16'b0000000000000010   ;
13'd431:weight<=16'b0000000000101110   ;
13'd432:weight<=16'b0000000000100100   ;
13'd433:weight<=16'b1111111101000011   ;
13'd434:weight<=16'b1111111111000100   ;
13'd435:weight<=16'b0000000001010011   ;
13'd436:weight<=16'b0000000011000101   ;
13'd437:weight<=16'b0000000011110010   ;
13'd438:weight<=16'b1111111110001010   ;
13'd439:weight<=16'b1111111101111011   ;
13'd440:weight<=16'b1111111101011100   ;
13'd441:weight<=16'b1111111111001101   ;
13'd442:weight<=16'b1111111111011101   ;
13'd443:weight<=16'b0000000001101010   ;
13'd444:weight<=16'b0000000001000110   ;
13'd445:weight<=16'b0000000010111011   ;
13'd446:weight<=16'b0000000000000000   ;
13'd447:weight<=16'b1111111111000001   ;
13'd448:weight<=16'b1111111110110000   ;
13'd449:weight<=16'b0000000000101111   ;
13'd450:weight<=16'b0000000010001100   ;
13'd451:weight<=16'b0000000001011111   ;
13'd452:weight<=16'b1111111111100101   ;
13'd453:weight<=16'b1111111111100100   ;
13'd454:weight<=16'b1111111111100001   ;
13'd455:weight<=16'b1111111110110111   ;
13'd456:weight<=16'b1111111110101110   ;
13'd457:weight<=16'b0000000000010010   ;
13'd458:weight<=16'b0000000001100010   ;
13'd459:weight<=16'b1111111110101011   ;
13'd460:weight<=16'b1111111111001001   ;
13'd461:weight<=16'b1111111110100011   ;
13'd462:weight<=16'b1111111110010011   ;
13'd463:weight<=16'b0000000010011011   ;
13'd464:weight<=16'b0000000000101001   ;
13'd465:weight<=16'b1111111111010011   ;
13'd466:weight<=16'b1111111111111101   ;
13'd467:weight<=16'b0000000011001100   ;
13'd468:weight<=16'b1111111111010011   ;
13'd469:weight<=16'b1111111111010001   ;
13'd470:weight<=16'b0000000010100010   ;
13'd471:weight<=16'b0000000001100001   ;
13'd472:weight<=16'b1111111101001011   ;
13'd473:weight<=16'b1111111111000010   ;
13'd474:weight<=16'b1111111101111111   ;
13'd475:weight<=16'b0000000001010000   ;
13'd476:weight<=16'b0000000000111010   ;
13'd477:weight<=16'b0000000100100000   ;
13'd478:weight<=16'b0000000000001000   ;
13'd479:weight<=16'b1111111101010010   ;
13'd480:weight<=16'b0000000001100000   ;
13'd481:weight<=16'b1111111111100110   ;
13'd482:weight<=16'b1111111111010101   ;
13'd483:weight<=16'b0000000110000101   ;
13'd484:weight<=16'b1111111101010011   ;
13'd485:weight<=16'b1111111110011001   ;
13'd486:weight<=16'b1111111111110111   ;
13'd487:weight<=16'b1111111111000110   ;
13'd488:weight<=16'b0000000000001101   ;
13'd489:weight<=16'b1111111111101011   ;
13'd490:weight<=16'b1111111101011100   ;
13'd491:weight<=16'b1111111111001101   ;
13'd492:weight<=16'b1111111111011101   ;
13'd493:weight<=16'b0000000001101010   ;
13'd494:weight<=16'b0000000001000110   ;
13'd495:weight<=16'b0000000010111011   ;
13'd496:weight<=16'b0000000000000000   ;
13'd497:weight<=16'b1111111111000001   ;
13'd498:weight<=16'b1111111110110000   ;
13'd499:weight<=16'b0000000000101111   ;
13'd500:weight<=16'b0000000000100110   ;
13'd501:weight<=16'b1111111110110001   ;
13'd502:weight<=16'b0000000011011011   ;
13'd503:weight<=16'b1111111110100001   ;
13'd504:weight<=16'b1111111111111000   ;
13'd505:weight<=16'b1111111111000011   ;
13'd506:weight<=16'b0000000010111100   ;
13'd507:weight<=16'b1111111111010011   ;
13'd508:weight<=16'b1111111111010001   ;
13'd509:weight<=16'b1111111110111100   ;
13'd510:weight<=16'b1111111111001001   ;
13'd511:weight<=16'b1111111110100011   ;
13'd512:weight<=16'b1111111110010011   ;
13'd513:weight<=16'b0000000010011011   ;
13'd514:weight<=16'b0000000000101001   ;
13'd515:weight<=16'b1111111111010011   ;
13'd516:weight<=16'b1111111111111101   ;
13'd517:weight<=16'b0000000011001100   ;
13'd518:weight<=16'b1111111111010011   ;
13'd519:weight<=16'b1111111111010001;
13'd520:weight<=16'b1111111110111010   ;
13'd521:weight<=16'b0000000001001111   ;
13'd522:weight<=16'b1111111100110101   ;
13'd523:weight<=16'b0000000101000011   ;
13'd524:weight<=16'b1111111101111101   ;
13'd525:weight<=16'b0000000000001101   ;
13'd526:weight<=16'b0000000000111111   ;
13'd527:weight<=16'b0000000011110110   ;
13'd528:weight<=16'b0000000001110000   ;
13'd529:weight<=16'b1111111010110011   ;
13'd530:weight<=16'b0000000001100000   ;
13'd531:weight<=16'b1111111111100110   ;
13'd532:weight<=16'b1111111111010101   ;
13'd533:weight<=16'b0000000110000101   ;
13'd534:weight<=16'b1111111101010011   ;
13'd535:weight<=16'b1111111110011001   ;
13'd536:weight<=16'b1111111111110111   ;
13'd537:weight<=16'b1111111111000110   ;
13'd538:weight<=16'b0000000000001101   ;
13'd539:weight<=16'b1111111111101011   ;
13'd540:weight<=16'b0000000000010001   ;
13'd541:weight<=16'b0000000000011110   ;
13'd542:weight<=16'b0000000000100100   ;
13'd543:weight<=16'b0000000001100100   ;
13'd544:weight<=16'b1111111110010110   ;
13'd545:weight<=16'b0000000000101101   ;
13'd546:weight<=16'b1111111111001100   ;
13'd547:weight<=16'b1111111110010001   ;
13'd548:weight<=16'b0000000001000011   ;
13'd549:weight<=16'b0000000000000110   ;
13'd550:weight<=16'b0000000000100110   ;
13'd551:weight<=16'b1111111110110001   ;
13'd552:weight<=16'b0000000011011011   ;
13'd553:weight<=16'b1111111110100001   ;
13'd554:weight<=16'b1111111111111000   ;
13'd555:weight<=16'b1111111111000011   ;
13'd556:weight<=16'b0000000010111100   ;
13'd557:weight<=16'b1111111111010011   ;
13'd558:weight<=16'b1111111111010001   ;
13'd559:weight<=16'b1111111110111100   ;
13'd560:weight<=16'b0000000010100011   ;
13'd561:weight<=16'b0000000000101111   ;
13'd562:weight<=16'b0000000001100001   ;
13'd563:weight<=16'b1111111110100111   ;
13'd564:weight<=16'b0000000000001110   ;
13'd565:weight<=16'b0000000000010111   ;
13'd566:weight<=16'b0000000001000110   ;
13'd567:weight<=16'b0000000000011001   ;
13'd568:weight<=16'b1111111010100101   ;
13'd569:weight<=16'b0000000000101101   ;
13'd570:weight<=16'b1111111110111010   ;
13'd571:weight<=16'b0000000001001111   ;
13'd572:weight<=16'b1111111100110101   ;
13'd573:weight<=16'b0000000101000011   ;
13'd574:weight<=16'b1111111101111101   ;
13'd575:weight<=16'b0000000000001101   ;
13'd576:weight<=16'b0000000000111111   ;
13'd577:weight<=16'b0000000011110110   ;
13'd578:weight<=16'b0000000001110000   ;
13'd579:weight<=16'b1111111010110011   ;
13'd580:weight<=16'b1111111110011011   ;
13'd581:weight<=16'b0000000001100101   ;
13'd582:weight<=16'b0000000101000001   ;
13'd583:weight<=16'b1111111101001011   ;
13'd584:weight<=16'b0000000001001101   ;
13'd585:weight<=16'b0000000001101100   ;
13'd586:weight<=16'b1111111111011100   ;
13'd587:weight<=16'b1111111101011111   ;
13'd588:weight<=16'b0000000000011000   ;
13'd589:weight<=16'b1111111110001001   ;
13'd590:weight<=16'b0000000000010001   ;
13'd591:weight<=16'b0000000000011110   ;
13'd592:weight<=16'b0000000000100100   ;
13'd593:weight<=16'b0000000001100100   ;
13'd594:weight<=16'b1111111110010110   ;
13'd595:weight<=16'b0000000000101101   ;
13'd596:weight<=16'b1111111111001100   ;
13'd597:weight<=16'b1111111110010001   ;
13'd598:weight<=16'b0000000001000011   ;
13'd599:weight<=16'b0000000000000110   ;
13'd600:weight<=16'b0000000000010000   ;
13'd601:weight<=16'b1111111111111110   ;
13'd602:weight<=16'b1111111110110000   ;
13'd603:weight<=16'b0000000001100101   ;
13'd604:weight<=16'b0000000000000000   ;
13'd605:weight<=16'b1111111111101010   ;
13'd606:weight<=16'b0000000001111011   ;
13'd607:weight<=16'b1111111110100001   ;
13'd608:weight<=16'b1111111111000100   ;
13'd609:weight<=16'b0000000000110101   ;
13'd610:weight<=16'b0000000010100011   ;
13'd611:weight<=16'b0000000000101111   ;
13'd612:weight<=16'b0000000001100001   ;
13'd613:weight<=16'b1111111110100111   ;
13'd614:weight<=16'b0000000000001110   ;
13'd615:weight<=16'b0000000000010111   ;
13'd616:weight<=16'b0000000001000110   ;
13'd617:weight<=16'b0000000000011001   ;
13'd618:weight<=16'b1111111010100101   ;
13'd619:weight<=16'b0000000000101101   ;
13'd620:weight<=16'b1111111110001000   ;
13'd621:weight<=16'b1111111101000111   ;
13'd622:weight<=16'b0000000000011010   ;
13'd623:weight<=16'b0000000000100100   ;
13'd624:weight<=16'b0000000001101100   ;
13'd625:weight<=16'b0000000010001011   ;
13'd626:weight<=16'b0000000001001000   ;
13'd627:weight<=16'b0000000001000001   ;
13'd628:weight<=16'b1111111101110111   ;
13'd629:weight<=16'b0000000000100011   ;
13'd630:weight<=16'b1111111110011011   ;
13'd631:weight<=16'b0000000001100101   ;
13'd632:weight<=16'b0000000101000001   ;
13'd633:weight<=16'b1111111101001011   ;
13'd634:weight<=16'b0000000001001101   ;
13'd635:weight<=16'b0000000001101100   ;
13'd636:weight<=16'b1111111111011100   ;
13'd637:weight<=16'b1111111101011111   ;
13'd638:weight<=16'b0000000000011000   ;
13'd639:weight<=16'b1111111110001001   ;
13'd640:weight<=16'b1111111101111111   ;
13'd641:weight<=16'b1111111011010100   ;
13'd642:weight<=16'b0000000000111110   ;
13'd643:weight<=16'b0000000011000101   ;
13'd644:weight<=16'b1111111110110010   ;
13'd645:weight<=16'b1111111111101101   ;
13'd646:weight<=16'b0000000010000101   ;
13'd647:weight<=16'b0000000001000111   ;
13'd648:weight<=16'b1111111111110100   ;
13'd649:weight<=16'b0000000001100001   ;
13'd650:weight<=16'b0000000000010000   ;
13'd651:weight<=16'b1111111111111110   ;
13'd652:weight<=16'b1111111110110000   ;
13'd653:weight<=16'b0000000001100101   ;
13'd654:weight<=16'b0000000000000000   ;
13'd655:weight<=16'b1111111111101010   ;
13'd656:weight<=16'b0000000001111011   ;
13'd657:weight<=16'b1111111110100001   ;
13'd658:weight<=16'b1111111111000100   ;
13'd659:weight<=16'b0000000000110101   ;
13'd660:weight<=16'b0000000000001000   ;
13'd661:weight<=16'b0000000000000101   ;
13'd662:weight<=16'b1111111110010100   ;
13'd663:weight<=16'b0000000000011010   ;
13'd664:weight<=16'b1111111111001011   ;
13'd665:weight<=16'b0000000001011111   ;
13'd666:weight<=16'b0000000000000111   ;
13'd667:weight<=16'b0000000010000010   ;
13'd668:weight<=16'b0000000001001111   ;
13'd669:weight<=16'b1111111101100100   ;
13'd670:weight<=16'b1111111110001000   ;
13'd671:weight<=16'b1111111101000111   ;
13'd672:weight<=16'b0000000000011010   ;
13'd673:weight<=16'b0000000000100100   ;
13'd674:weight<=16'b0000000001101100   ;
13'd675:weight<=16'b0000000010001011   ;
13'd676:weight<=16'b0000000001001000   ;
13'd677:weight<=16'b0000000001000001   ;
13'd678:weight<=16'b1111111101110111   ;
13'd679:weight<=16'b0000000000100011   ;
13'd680:weight<=16'b1111111110110110   ;
13'd681:weight<=16'b0000000010001110   ;
13'd682:weight<=16'b0000000001110101   ;
13'd683:weight<=16'b1111111110001101   ;
13'd684:weight<=16'b0000000001000011   ;
13'd685:weight<=16'b1111111110011001   ;
13'd686:weight<=16'b1111111111011100   ;
13'd687:weight<=16'b1111111101111011   ;
13'd688:weight<=16'b0000000001110110   ;
13'd689:weight<=16'b0000000000111001   ;
13'd690:weight<=16'b1111111101111111   ;
13'd691:weight<=16'b1111111011010100   ;
13'd692:weight<=16'b0000000000111110   ;
13'd693:weight<=16'b0000000011000101   ;
13'd694:weight<=16'b1111111110110010   ;
13'd695:weight<=16'b1111111111101101   ;
13'd696:weight<=16'b0000000010000101   ;
13'd697:weight<=16'b0000000001000111   ;
13'd698:weight<=16'b1111111111110100   ;
13'd699:weight<=16'b0000000001100001   ;
13'd700:weight<=16'b1111111110010010   ;
13'd701:weight<=16'b1111111111110111   ;
13'd702:weight<=16'b0000000010000000   ;
13'd703:weight<=16'b0000000000001011   ;
13'd704:weight<=16'b0000000010000100   ;
13'd705:weight<=16'b1111111111111011   ;
13'd706:weight<=16'b0000000000000011   ;
13'd707:weight<=16'b1111111110001100   ;
13'd708:weight<=16'b1111111110111001   ;
13'd709:weight<=16'b0000000000110010   ;
13'd710:weight<=16'b0000000000001000   ;
13'd711:weight<=16'b0000000000000101   ;
13'd712:weight<=16'b1111111110010100   ;
13'd713:weight<=16'b0000000000011010   ;
13'd714:weight<=16'b1111111111001011   ;
13'd715:weight<=16'b0000000001011111   ;
13'd716:weight<=16'b0000000000000111   ;
13'd717:weight<=16'b0000000010000010   ;
13'd718:weight<=16'b0000000001001111   ;
13'd719:weight<=16'b1111111101100100   ;
13'd720:weight<=16'b1111111111011111   ;
13'd721:weight<=16'b1111111110100010   ;
13'd722:weight<=16'b0000000001011111   ;
13'd723:weight<=16'b1111111011011101   ;
13'd724:weight<=16'b1111111110110000   ;
13'd725:weight<=16'b0000000011101001   ;
13'd726:weight<=16'b0000000101010100   ;
13'd727:weight<=16'b0000000000000010   ;
13'd728:weight<=16'b0000000010001111   ;
13'd729:weight<=16'b1111111011001101   ;
13'd730:weight<=16'b1111111110110110   ;
13'd731:weight<=16'b0000000010001110   ;
13'd732:weight<=16'b0000000001110101   ;
13'd733:weight<=16'b1111111110001101   ;
13'd734:weight<=16'b0000000001000011   ;
13'd735:weight<=16'b1111111110011001   ;
13'd736:weight<=16'b1111111111011100   ;
13'd737:weight<=16'b1111111101111011   ;
13'd738:weight<=16'b0000000001110110   ;
13'd739:weight<=16'b0000000000111001   ;
13'd740:weight<=16'b0000000001110011   ;
13'd741:weight<=16'b1111111101000000   ;
13'd742:weight<=16'b1111111110100111   ;
13'd743:weight<=16'b0000000001011011   ;
13'd744:weight<=16'b0000000001101110   ;
13'd745:weight<=16'b0000000000110101   ;
13'd746:weight<=16'b1111111111011100   ;
13'd747:weight<=16'b1111111111010010   ;
13'd748:weight<=16'b1111111110001011   ;
13'd749:weight<=16'b0000000001110100   ;
13'd750:weight<=16'b1111111110010010   ;
13'd751:weight<=16'b1111111111110111   ;
13'd752:weight<=16'b0000000010000000   ;
13'd753:weight<=16'b0000000000001011   ;
13'd754:weight<=16'b0000000010000100   ;
13'd755:weight<=16'b1111111111111011   ;
13'd756:weight<=16'b0000000000000011   ;
13'd757:weight<=16'b1111111110001100   ;
13'd758:weight<=16'b1111111110111001   ;
13'd759:weight<=16'b0000000000110010   ;
13'd760:weight<=16'b1111111110001111   ;
13'd761:weight<=16'b0000000001011111   ;
13'd762:weight<=16'b0000000001000001   ;
13'd763:weight<=16'b0000000001111000   ;
13'd764:weight<=16'b0000000000011110   ;
13'd765:weight<=16'b0000000001110110   ;
13'd766:weight<=16'b0000000000010100   ;
13'd767:weight<=16'b1111111111100110   ;
13'd768:weight<=16'b1111111110100101   ;
13'd769:weight<=16'b1111111101001011   ;
13'd770:weight<=16'b1111111111011111   ;
13'd771:weight<=16'b1111111110100010   ;
13'd772:weight<=16'b0000000001011111   ;
13'd773:weight<=16'b1111111011011101   ;
13'd774:weight<=16'b1111111110110000   ;
13'd775:weight<=16'b0000000011101001   ;
13'd776:weight<=16'b0000000101010100   ;
13'd777:weight<=16'b0000000000000010   ;
13'd778:weight<=16'b0000000010001111   ;
13'd779:weight<=16'b1111111011001101   ;
13'd780:weight<=16'b1111111110110010   ;
13'd781:weight<=16'b1111111110011000   ;
13'd782:weight<=16'b1111111110010001   ;
13'd783:weight<=16'b0000000011111101   ;
13'd784:weight<=16'b0000001000100011   ;
13'd785:weight<=16'b1111111101000001   ;
13'd786:weight<=16'b0000000001001000   ;
13'd787:weight<=16'b1111111101100001   ;
13'd788:weight<=16'b1111111101100010   ;
13'd789:weight<=16'b1111111111110101   ;
13'd790:weight<=16'b0000000001110011   ;
13'd791:weight<=16'b1111111101000000   ;
13'd792:weight<=16'b1111111110100111   ;
13'd793:weight<=16'b0000000001011011   ;
13'd794:weight<=16'b0000000001101110   ;
13'd795:weight<=16'b0000000000110101   ;
13'd796:weight<=16'b1111111111011100   ;
13'd797:weight<=16'b1111111111010010   ;
13'd798:weight<=16'b1111111110001011   ;
13'd799:weight<=16'b0000000001110100   ;
13'd800:weight<=16'b0000000001001001   ;
13'd801:weight<=16'b0000000000001101   ;
13'd802:weight<=16'b1111111111110011   ;
13'd803:weight<=16'b0000000001101001   ;
13'd804:weight<=16'b1111111110111001   ;
13'd805:weight<=16'b1111111101010011   ;
13'd806:weight<=16'b0000000001011011   ;
13'd807:weight<=16'b0000000000011111   ;
13'd808:weight<=16'b1111111101110000   ;
13'd809:weight<=16'b0000000010010000   ;
13'd810:weight<=16'b1111111110001111   ;
13'd811:weight<=16'b0000000001011111   ;
13'd812:weight<=16'b0000000001000001   ;
13'd813:weight<=16'b0000000001111000   ;
13'd814:weight<=16'b0000000000011110   ;
13'd815:weight<=16'b0000000001110110   ;
13'd816:weight<=16'b0000000000010100   ;
13'd817:weight<=16'b1111111111100110   ;
13'd818:weight<=16'b1111111110100101   ;
13'd819:weight<=16'b1111111101001011   ;
13'd820:weight<=16'b0000000000010100   ;
13'd821:weight<=16'b1111111101001100   ;
13'd822:weight<=16'b0000000010110111   ;
13'd823:weight<=16'b1111111111001010   ;
13'd824:weight<=16'b0000000011111110   ;
13'd825:weight<=16'b0000000000001110   ;
13'd826:weight<=16'b1111111010100001   ;
13'd827:weight<=16'b1111111111010011   ;
13'd828:weight<=16'b1111111110110011   ;
13'd829:weight<=16'b0000000011001101   ;
13'd830:weight<=16'b1111111110110010   ;
13'd831:weight<=16'b1111111110011000   ;
13'd832:weight<=16'b1111111110010001  ;
13'd833:weight<=16'b0000000011111101   ;
13'd834:weight<=16'b0000001000100011   ;
13'd835:weight<=16'b1111111101000001   ;
13'd836:weight<=16'b0000000001001000   ;
13'd837:weight<=16'b1111111101100001   ;
13'd838:weight<=16'b1111111101100010   ;
13'd839:weight<=16'b1111111111110101   ;
13'd840:weight<=16'b0000000000110101   ;
13'd841:weight<=16'b1111111101011100   ;
13'd842:weight<=16'b1111111111110111   ;
13'd843:weight<=16'b0000000000000000   ;
13'd844:weight<=16'b0000000010011001   ;
13'd845:weight<=16'b1111111111101111   ;
13'd846:weight<=16'b1111111101010000   ;
13'd847:weight<=16'b0000000000010101   ;
13'd848:weight<=16'b0000000000000001   ;
13'd849:weight<=16'b0000000010000111   ;
13'd850:weight<=16'b0000000001001001   ;
13'd851:weight<=16'b0000000000001101   ;
13'd852:weight<=16'b1111111111110011   ;
13'd853:weight<=16'b0000000001101001   ;
13'd854:weight<=16'b1111111110111001   ;
13'd855:weight<=16'b1111111101010011   ;
13'd856:weight<=16'b0000000001011011   ;
13'd857:weight<=16'b0000000000011111   ;
13'd858:weight<=16'b1111111101110000  ;
13'd859:weight<=16'b0000000010010000   ;
13'd860:weight<=16'b0000000000100001   ;
13'd861:weight<=16'b0000000100011100   ;
13'd862:weight<=16'b1111111111100010   ;
13'd863:weight<=16'b1111111111110110   ;
13'd864:weight<=16'b1111111110100001   ;
13'd865:weight<=16'b0000000001010111   ;
13'd866:weight<=16'b1111111110000000   ;
13'd867:weight<=16'b0000000000100100   ;
13'd868:weight<=16'b1111111111100111   ;
13'd869:weight<=16'b1111111110010001   ;
13'd870:weight<=16'b0000000000010100   ;
13'd871:weight<=16'b1111111101001100   ;
13'd872:weight<=16'b0000000010110111   ;
13'd873:weight<=16'b1111111111001010   ;
13'd874:weight<=16'b0000000011111110   ;
13'd875:weight<=16'b0000000000001110   ;
13'd876:weight<=16'b1111111010100001   ;
13'd877:weight<=16'b1111111111010011   ;
13'd878:weight<=16'b1111111110110011   ;
13'd879:weight<=16'b0000000011001101   ;
13'd880:weight<=16'b1111111111011111   ;
13'd881:weight<=16'b1111111111111100   ;
13'd882:weight<=16'b0000000001010111   ;
13'd883:weight<=16'b0000000000110000   ;
13'd884:weight<=16'b1111111111000101   ;
13'd885:weight<=16'b1111111111010011   ;
13'd886:weight<=16'b1111111110110111   ;
13'd887:weight<=16'b0000000010010111   ;
13'd888:weight<=16'b0000000001011110   ;
13'd889:weight<=16'b1111111101111010   ;
13'd890:weight<=16'b0000000000110101   ;
13'd891:weight<=16'b1111111101011100   ;
13'd892:weight<=16'b1111111111110111   ;
13'd893:weight<=16'b0000000000000000   ;
13'd894:weight<=16'b0000000010011001   ;
13'd895:weight<=16'b1111111111101111   ;
13'd896:weight<=16'b1111111101010000   ;
13'd897:weight<=16'b0000000000010101   ;
13'd898:weight<=16'b0000000000000001   ;
13'd899:weight<=16'b0000000010000111   ;
13'd900:weight<=16'b1111111111010000   ;
13'd901:weight<=16'b0000000010000101   ;
13'd902:weight<=16'b1111111110110101   ;
13'd903:weight<=16'b0000000010001101   ;
13'd904:weight<=16'b1111111110000001   ;
13'd905:weight<=16'b1111111110101101   ;
13'd906:weight<=16'b0000000010100111   ;
13'd907:weight<=16'b1111111111011111   ;
13'd908:weight<=16'b1111111100100100   ;
13'd909:weight<=16'b0000000010111110   ;
13'd910:weight<=16'b0000000000100001   ;
13'd911:weight<=16'b0000000100011100   ;
13'd912:weight<=16'b1111111111100010   ;
13'd913:weight<=16'b1111111111110110   ;
13'd914:weight<=16'b1111111110100001   ;
13'd915:weight<=16'b0000000001010111   ;
13'd916:weight<=16'b1111111110000000   ;
13'd917:weight<=16'b0000000000100100   ;
13'd918:weight<=16'b1111111111100111   ;
13'd919:weight<=16'b1111111110010001   ;
13'd920:weight<=16'b0000000000000000   ;
13'd921:weight<=16'b1111111110101001   ;
13'd922:weight<=16'b0000000011010111   ;
13'd923:weight<=16'b1111111101110010   ;
13'd924:weight<=16'b1111111110011101   ;
13'd925:weight<=16'b1111111110001011   ;
13'd926:weight<=16'b0000000010011001   ;
13'd927:weight<=16'b1111111111010010   ;
13'd928:weight<=16'b1111111101000110   ;
13'd929:weight<=16'b0000000101000010   ;
13'd930:weight<=16'b1111111111011111   ;
13'd931:weight<=16'b1111111111111100   ;
13'd932:weight<=16'b0000000001010111   ;
13'd933:weight<=16'b0000000000110000   ;
13'd934:weight<=16'b1111111111000101   ;
13'd935:weight<=16'b1111111111010011   ;
13'd936:weight<=16'b1111111110110111   ;
13'd937:weight<=16'b0000000010010111   ;
13'd938:weight<=16'b0000000001011110   ;
13'd939:weight<=16'b1111111101111010   ;
13'd940:weight<=16'b0000000011011100   ;
13'd941:weight<=16'b1111111100111110   ;
13'd942:weight<=16'b1111111001000000   ;
13'd943:weight<=16'b0000001000000011   ;
13'd944:weight<=16'b1111111101100101   ;
13'd945:weight<=16'b1111111010001100   ;
13'd946:weight<=16'b1111111110111011   ;
13'd947:weight<=16'b0000001001000011   ;
13'd948:weight<=16'b0000000011010101   ;
13'd949:weight<=16'b1111111101110000   ;
13'd950:weight<=16'b1111111111010000   ;
13'd951:weight<=16'b0000000010000101   ;
13'd952:weight<=16'b1111111110110101   ;
13'd953:weight<=16'b0000000010001101   ;
13'd954:weight<=16'b1111111110000001   ;
13'd955:weight<=16'b1111111110101101   ;
13'd956:weight<=16'b0000000010100111   ;
13'd957:weight<=16'b1111111111011111   ;
13'd958:weight<=16'b1111111100100100   ;
13'd959:weight<=16'b0000000010111110   ;
13'd960:weight<=16'b1111111111010010   ;
13'd961:weight<=16'b0000000000010100   ;
13'd962:weight<=16'b1111111111110101   ;
13'd963:weight<=16'b0000000000111101   ;
13'd964:weight<=16'b1111111110001111   ;
13'd965:weight<=16'b1111111101010011   ;
13'd966:weight<=16'b0000000001011100   ;
13'd967:weight<=16'b0000000000101111   ;
13'd968:weight<=16'b0000000010100100   ;
13'd969:weight<=16'b1111111111011111   ;
13'd970:weight<=16'b0000000000000000   ;
13'd971:weight<=16'b1111111110101001   ;
13'd972:weight<=16'b0000000011010111   ;
13'd973:weight<=16'b1111111101110010   ;
13'd974:weight<=16'b1111111110011101   ;
13'd975:weight<=16'b1111111110001011   ;
13'd976:weight<=16'b0000000010011001   ;
13'd977:weight<=16'b1111111111010010   ;
13'd978:weight<=16'b1111111101000110   ;
13'd979:weight<=16'b0000000101000010   ;
13'd980:weight<=16'b1111111111000110   ;
13'd981:weight<=16'b0000000001101101   ;
13'd982:weight<=16'b1111111101011010   ;
13'd983:weight<=16'b0000000001010111   ;
13'd984:weight<=16'b1111111111101001   ;
13'd985:weight<=16'b0000000001111110   ;
13'd986:weight<=16'b0000000010111100   ;
13'd987:weight<=16'b1111111111101111   ;
13'd988:weight<=16'b1111111111001111   ;
13'd989:weight<=16'b1111111110100100   ;
13'd990:weight<=16'b0000000011011100   ;
13'd991:weight<=16'b1111111100111110   ;
13'd992:weight<=16'b1111111001000000   ;
13'd993:weight<=16'b0000001000000011   ;
13'd994:weight<=16'b1111111101100101   ;
13'd995:weight<=16'b1111111010001100   ;
13'd996:weight<=16'b1111111110111011   ;
13'd997:weight<=16'b0000001001000011   ;
13'd998:weight<=16'b0000000011010101   ;
13'd999:weight<=16'b1111111101110000   ;
13'd1000:weight<=16'b0000000000100110   ;
13'd1001:weight<=16'b0000000001100010   ;
13'd1002:weight<=16'b1111111101110000   ;
13'd1003:weight<=16'b0000000011001011   ;
13'd1004:weight<=16'b1111111111010011   ;
13'd1005:weight<=16'b1111111111101011  ;
13'd1006:weight<=16'b0000000000000011   ;
13'd1007:weight<=16'b0000000001011010   ;
13'd1008:weight<=16'b1111111110000101   ;
13'd1009:weight<=16'b1111111110111101   ;
13'd1010:weight<=16'b1111111111010010   ;
13'd1011:weight<=16'b0000000000010100   ;
13'd1012:weight<=16'b1111111111110101   ;
13'd1013:weight<=16'b0000000000111101   ;
13'd1014:weight<=16'b1111111110001111   ;
13'd1015:weight<=16'b1111111101010011   ;
13'd1016:weight<=16'b0000000001011100   ;
13'd1017:weight<=16'b0000000000101111   ;
13'd1018:weight<=16'b0000000010100100   ;
13'd1019:weight<=16'b1111111111011111   ;
13'd1020:weight<=16'b0000000001000011   ;
13'd1021:weight<=16'b0000000100000001   ;
13'd1022:weight<=16'b1111111100001001   ;
13'd1023:weight<=16'b1111111111010111   ;
13'd1024:weight<=16'b1111111100001010   ;
13'd1025:weight<=16'b1111111100001011   ;
13'd1026:weight<=16'b0000000100001010   ;
13'd1027:weight<=16'b0000000100111100   ;
13'd1028:weight<=16'b1111111101101100   ;
13'd1029:weight<=16'b0000000001100001   ;
13'd1030:weight<=16'b1111111111000110   ;
13'd1031:weight<=16'b0000000001101101   ;
13'd1032:weight<=16'b1111111101011010   ;
13'd1033:weight<=16'b0000000001010111   ;
13'd1034:weight<=16'b1111111111101001   ;
13'd1035:weight<=16'b0000000001111110   ;
13'd1036:weight<=16'b0000000010111100   ;
13'd1037:weight<=16'b1111111111101111   ;
13'd1038:weight<=16'b1111111111001111   ;
13'd1039:weight<=16'b1111111110100100   ;
13'd1040:weight<=16'b1111111010100100   ;
13'd1041:weight<=16'b1111111101111110   ;
13'd1042:weight<=16'b0000000000000100   ;
13'd1043:weight<=16'b1111111101110000   ;
13'd1044:weight<=16'b0000000000101100   ;
13'd1045:weight<=16'b0000000100000011   ;
13'd1046:weight<=16'b1111111111100010   ;
13'd1047:weight<=16'b1111111111011110   ;
13'd1048:weight<=16'b0000000000110001   ;
13'd1049:weight<=16'b0000000101110100   ;
13'd1050:weight<=16'b0000000000100110   ;
13'd1051:weight<=16'b0000000001100010   ;
13'd1052:weight<=16'b1111111101110000   ;
13'd1053:weight<=16'b0000000011001011   ;
13'd1054:weight<=16'b1111111111010011   ;
13'd1055:weight<=16'b1111111111101011   ;
13'd1056:weight<=16'b0000000000000011   ;
13'd1057:weight<=16'b0000000001011010   ;
13'd1058:weight<=16'b1111111110000101   ;
13'd1059:weight<=16'b1111111110111101   ;
13'd1060:weight<=16'b1111111111000100   ;
13'd1061:weight<=16'b0000000010101010   ;
13'd1062:weight<=16'b0000000000000001   ;
13'd1063:weight<=16'b1111111110010011   ;
13'd1064:weight<=16'b0000000000001101   ;
13'd1065:weight<=16'b0000000010000010   ;
13'd1066:weight<=16'b1111111111110010   ;
13'd1067:weight<=16'b0000000001101010   ;
13'd1068:weight<=16'b1111111101100101   ;
13'd1069:weight<=16'b0000000000010011   ;
13'd1070:weight<=16'b0000000001000011   ;
13'd1071:weight<=16'b0000000100000001   ;
13'd1072:weight<=16'b1111111100001001   ;
13'd1073:weight<=16'b1111111111010111   ;
13'd1074:weight<=16'b1111111100001010   ;
13'd1075:weight<=16'b1111111100001011   ;
13'd1076:weight<=16'b0000000100001010   ;
13'd1077:weight<=16'b0000000100111100   ;
13'd1078:weight<=16'b1111111101101100   ;
13'd1079:weight<=16'b0000000001100001   ;
13'd1080:weight<=16'b1111111111000101   ;
13'd1081:weight<=16'b0000000000010001   ;
13'd1082:weight<=16'b1111111111010100   ;
13'd1083:weight<=16'b1111111111101011   ;
13'd1084:weight<=16'b0000000000011001   ;
13'd1085:weight<=16'b0000000001011101   ;
13'd1086:weight<=16'b0000000001000011   ;
13'd1087:weight<=16'b1111111111011010   ;
13'd1088:weight<=16'b1111111101110110   ;
13'd1089:weight<=16'b0000000001111110   ;
13'd1090:weight<=16'b1111111010100100   ;
13'd1091:weight<=16'b1111111101111110   ;
13'd1092:weight<=16'b0000000000000100   ;
13'd1093:weight<=16'b1111111101110000   ;
13'd1094:weight<=16'b0000000000101100   ;
13'd1095:weight<=16'b0000000100000011   ;
13'd1096:weight<=16'b1111111111100010   ;
13'd1097:weight<=16'b1111111111011110   ;
13'd1098:weight<=16'b0000000000110001   ;
13'd1099:weight<=16'b0000000101110100   ;
13'd1100:weight<=16'b1111111111010010   ;
13'd1101:weight<=16'b1111111110111000   ;
13'd1102:weight<=16'b0000000001101101   ;
13'd1103:weight<=16'b1111111100011010   ;
13'd1104:weight<=16'b0000000010010110   ;
13'd1105:weight<=16'b0000000101100011   ;
13'd1106:weight<=16'b1111111101101000   ;
13'd1107:weight<=16'b0000000010011101   ;
13'd1108:weight<=16'b1111111101100111   ;
13'd1109:weight<=16'b1111111111001100   ;
13'd1110:weight<=16'b1111111111000100   ;
13'd1111:weight<=16'b0000000010101010   ;
13'd1112:weight<=16'b0000000000000001   ;
13'd1113:weight<=16'b1111111110010011   ;
13'd1114:weight<=16'b0000000000001101   ;
13'd1115:weight<=16'b0000000010000010   ;
13'd1116:weight<=16'b1111111111110010   ;
13'd1117:weight<=16'b0000000001101010   ;
13'd1118:weight<=16'b1111111101100101   ;
13'd1119:weight<=16'b0000000000010011   ;
13'd1120:weight<=16'b1111111110011101   ;
13'd1121:weight<=16'b1111111111011001   ;
13'd1122:weight<=16'b0000000001111101   ;
13'd1123:weight<=16'b1111111111111100   ;
13'd1124:weight<=16'b0000000001010110   ;
13'd1125:weight<=16'b1111111111010110   ;
13'd1126:weight<=16'b0000000000110101   ;
13'd1127:weight<=16'b1111111110110010   ;
13'd1128:weight<=16'b1111111110111111   ;
13'd1129:weight<=16'b0000000010100101   ;
13'd1130:weight<=16'b1111111111000101   ;
13'd1131:weight<=16'b0000000000010001   ;
13'd1132:weight<=16'b1111111111010100   ;
13'd1133:weight<=16'b1111111111101011   ;
13'd1134:weight<=16'b0000000000011001   ;
13'd1135:weight<=16'b0000000001011101   ;
13'd1136:weight<=16'b0000000001000011   ;
13'd1137:weight<=16'b1111111111011010   ;
13'd1138:weight<=16'b1111111101110110   ;
13'd1139:weight<=16'b0000000001111110   ;
13'd1140:weight<=16'b0000000001000010   ;
13'd1141:weight<=16'b0000000010001001   ;
13'd1142:weight<=16'b1111111111110111   ;
13'd1143:weight<=16'b0000000000000100   ;
13'd1144:weight<=16'b1111111110111100   ;
13'd1145:weight<=16'b1111111101110100   ;
13'd1146:weight<=16'b0000000011100010   ;
13'd1147:weight<=16'b1111111110000011   ;
13'd1148:weight<=16'b1111111111010010   ;
13'd1149:weight<=16'b1111111111110101   ;
13'd1150:weight<=16'b1111111111010010   ;
13'd1151:weight<=16'b1111111110111000   ;
13'd1152:weight<=16'b0000000001101101   ;
13'd1153:weight<=16'b1111111100011010   ;
13'd1154:weight<=16'b0000000010010110   ;
13'd1155:weight<=16'b0000000101100011   ;
13'd1156:weight<=16'b1111111101101000   ;
13'd1157:weight<=16'b0000000010011101   ;
13'd1158:weight<=16'b1111111101100111   ;
13'd1159:weight<=16'b1111111111001100   ;
13'd1160:weight<=16'b0000000000010011   ;
13'd1161:weight<=16'b0000000011101011   ;
13'd1162:weight<=16'b1111111011000100   ;
13'd1163:weight<=16'b0000000010100001   ;
13'd1164:weight<=16'b1111111010111001   ;
13'd1165:weight<=16'b1111111100011011   ;
13'd1166:weight<=16'b0000000101110010   ;
13'd1167:weight<=16'b0000000010001011   ;
13'd1168:weight<=16'b1111111101000000   ;
13'd1169:weight<=16'b0000000011010100   ;
13'd1170:weight<=16'b1111111110011101   ;
13'd1171:weight<=16'b1111111111011001   ;
13'd1172:weight<=16'b0000000001111101   ;
13'd1173:weight<=16'b1111111111111100   ;
13'd1174:weight<=16'b0000000001010110   ;
13'd1175:weight<=16'b1111111111010110   ;
13'd1176:weight<=16'b0000000000110101   ;
13'd1177:weight<=16'b1111111110110010   ;
13'd1178:weight<=16'b1111111110111111   ;
13'd1179:weight<=16'b0000000010100101   ;
13'd1180:weight<=16'b0000000000110001   ;
13'd1181:weight<=16'b1111111111101100   ;
13'd1182:weight<=16'b1111111111011101   ;
13'd1183:weight<=16'b0000000001101101   ;
13'd1184:weight<=16'b1111111110000011   ;
13'd1185:weight<=16'b0000000000001000   ;
13'd1186:weight<=16'b0000000001101101   ;
13'd1187:weight<=16'b0000000010000000   ;
13'd1188:weight<=16'b1111111111100111   ;
13'd1189:weight<=16'b1111111110000000   ;
13'd1190:weight<=16'b0000000001000010   ;
13'd1191:weight<=16'b0000000010001001   ;
13'd1192:weight<=16'b1111111111110111   ;
13'd1193:weight<=16'b0000000000000100   ;
13'd1194:weight<=16'b1111111110111100   ;
13'd1195:weight<=16'b1111111101110100   ;
13'd1196:weight<=16'b0000000011100010   ;
13'd1197:weight<=16'b1111111110000011   ;
13'd1198:weight<=16'b1111111111010010   ;
13'd1199:weight<=16'b1111111111110101   ;
13'd1200:weight<=16'b0000000010000001   ;
13'd1201:weight<=16'b0000000000000111   ;
13'd1202:weight<=16'b0000000000100000   ;
13'd1203:weight<=16'b1111111111001000   ;
13'd1204:weight<=16'b0000000000100111   ;
13'd1205:weight<=16'b1111111110010110   ;
13'd1206:weight<=16'b0000000010011100   ;
13'd1207:weight<=16'b1111111110001101   ;
13'd1208:weight<=16'b1111111111010011   ;
13'd1209:weight<=16'b1111111111101101   ;
13'd1210:weight<=16'b0000000000010011   ;
13'd1211:weight<=16'b0000000011101011   ;
13'd1212:weight<=16'b1111111011000100   ;
13'd1213:weight<=16'b0000000010100001   ;
13'd1214:weight<=16'b1111111010111001   ;
13'd1215:weight<=16'b1111111100011011   ;
13'd1216:weight<=16'b0000000101110010   ;
13'd1217:weight<=16'b0000000010001011   ;
13'd1218:weight<=16'b1111111101000000   ;
13'd1219:weight<=16'b0000000011010100   ;
13'd1220:weight<=16'b0000000000000100   ;
13'd1221:weight<=16'b1111111101100000   ;
13'd1222:weight<=16'b0000000000010101   ;
13'd1223:weight<=16'b1111111011000110   ;
13'd1224:weight<=16'b1111111111001000   ;
13'd1225:weight<=16'b0000000011101010   ;
13'd1226:weight<=16'b1111111111100111   ;
13'd1227:weight<=16'b0000000101001100   ;
13'd1228:weight<=16'b1111111111000110   ;
13'd1229:weight<=16'b0000000000110001   ;
13'd1230:weight<=16'b0000000000110001   ;
13'd1231:weight<=16'b1111111111101100   ;
13'd1232:weight<=16'b1111111111011101   ;
13'd1233:weight<=16'b0000000001101101   ;
13'd1234:weight<=16'b1111111110000011   ;
13'd1235:weight<=16'b0000000000001000   ;
13'd1236:weight<=16'b0000000001101101   ;
13'd1237:weight<=16'b0000000010000000   ;
13'd1238:weight<=16'b1111111111100111   ;
13'd1239:weight<=16'b1111111110000000   ;
13'd1240:weight<=16'b1111111111010001   ;
13'd1241:weight<=16'b0000000001010110   ;
13'd1242:weight<=16'b1111111111110111   ;
13'd1243:weight<=16'b1111111110010011   ;
13'd1244:weight<=16'b0000000001010000   ;
13'd1245:weight<=16'b1111111111011110   ;
13'd1246:weight<=16'b0000000001001000   ;
13'd1247:weight<=16'b1111111111010010   ;
13'd1248:weight<=16'b1111111111011010   ;
13'd1249:weight<=16'b0000000001010110   ;
13'd1250:weight<=16'b0000000010000001   ;
13'd1251:weight<=16'b0000000000000111   ;
13'd1252:weight<=16'b0000000000100000   ;
13'd1253:weight<=16'b1111111111001000   ;
13'd1254:weight<=16'b0000000000100111   ;
13'd1255:weight<=16'b1111111110010110   ;
13'd1256:weight<=16'b0000000010011100   ;
13'd1257:weight<=16'b1111111110001101   ;
13'd1258:weight<=16'b1111111111010011   ;
13'd1259:weight<=16'b1111111111101101   ;
13'd1260:weight<=16'b1111111111100011   ;
13'd1261:weight<=16'b0000000010100000   ;
13'd1262:weight<=16'b1111111111000000   ;
13'd1263:weight<=16'b1111111110101001   ;
13'd1264:weight<=16'b0000000000001000   ;
13'd1265:weight<=16'b1111111111110011   ;
13'd1266:weight<=16'b0000000000111101   ;
13'd1267:weight<=16'b0000000000100001   ;
13'd1268:weight<=16'b1111111111000000   ;
13'd1269:weight<=16'b0000000001100100   ;
13'd1270:weight<=16'b0000000000000100   ;
13'd1271:weight<=16'b1111111101100000   ;
13'd1272:weight<=16'b0000000000010101   ;
13'd1273:weight<=16'b1111111011000110   ;
13'd1274:weight<=16'b1111111111001000   ;
13'd1275:weight<=16'b0000000011101010   ;
13'd1276:weight<=16'b1111111111100111   ;
13'd1277:weight<=16'b0000000101001100   ;
13'd1278:weight<=16'b1111111111000110   ;
13'd1279:weight<=16'b0000000000110001   ;
13'd1280:weight<=16'b0000000011000110   ;
13'd1281:weight<=16'b1111111111001100   ;
13'd1282:weight<=16'b0000000000011111   ;
13'd1283:weight<=16'b0000000011011000   ;
13'd1284:weight<=16'b1111111111001001   ;
13'd1285:weight<=16'b1111111100101010   ;
13'd1286:weight<=16'b0000000000101100   ;
13'd1287:weight<=16'b1111111111010000   ;
13'd1288:weight<=16'b0000000000010001   ;
13'd1289:weight<=16'b1111111110110010   ;
13'd1290:weight<=16'b1111111111010001   ;
13'd1291:weight<=16'b0000000001010110   ;
13'd1292:weight<=16'b1111111111110111   ;
13'd1293:weight<=16'b1111111110010011   ;
13'd1294:weight<=16'b0000000001010000   ;
13'd1295:weight<=16'b1111111111011110   ;
13'd1296:weight<=16'b0000000001001000   ;
13'd1297:weight<=16'b1111111111010010   ;
13'd1298:weight<=16'b1111111111011010   ;
13'd1299:weight<=16'b0000000001010110   ;
13'd1300:weight<=16'b1111111100101011   ;
13'd1301:weight<=16'b0000010000011010   ;
13'd1302:weight<=16'b1111111110110010   ;
13'd1303:weight<=16'b1111111010110011   ;
13'd1304:weight<=16'b1111111100000000   ;
13'd1305:weight<=16'b0000000011101110   ;
13'd1306:weight<=16'b1111111101100001  ;
13'd1307:weight<=16'b1111111100110110   ;
13'd1308:weight<=16'b0000000001111101   ;
13'd1309:weight<=16'b0000000001001110   ;
13'd1310:weight<=16'b1111111111100011   ;
13'd1311:weight<=16'b0000000010100000   ;
13'd1312:weight<=16'b1111111111000000   ;
13'd1313:weight<=16'b1111111110101001   ;
13'd1314:weight<=16'b0000000000001000   ;
13'd1315:weight<=16'b1111111111110011   ;
13'd1316:weight<=16'b0000000000111101   ;
13'd1317:weight<=16'b0000000000100001   ;
13'd1318:weight<=16'b1111111111000000   ;
13'd1319:weight<=16'b0000000001100100   ;
13'd1320:weight<=16'b0000000001001011   ;
13'd1321:weight<=16'b0000000000000111   ;
13'd1322:weight<=16'b1111111111101110   ;
13'd1323:weight<=16'b1111111111111111   ;
13'd1324:weight<=16'b1111111111011000   ;
13'd1325:weight<=16'b1111111111111111   ;
13'd1326:weight<=16'b1111111111001110   ;
13'd1327:weight<=16'b0000000000111010   ;
13'd1328:weight<=16'b0000000001100000   ;
13'd1329:weight<=16'b1111111110110000   ;
13'd1330:weight<=16'b0000000011000110   ;
13'd1331:weight<=16'b1111111111001100   ;
13'd1332:weight<=16'b0000000000011111   ;
13'd1333:weight<=16'b0000000011011000   ;
13'd1334:weight<=16'b1111111111001001   ;
13'd1335:weight<=16'b1111111100101010   ;
13'd1336:weight<=16'b0000000000101100   ;
13'd1337:weight<=16'b1111111111010000   ;
13'd1338:weight<=16'b0000000000010001   ;
13'd1339:weight<=16'b1111111110110010   ;
13'd1340:weight<=16'b0000000011100111   ;
13'd1341:weight<=16'b1111111101111010   ;
13'd1342:weight<=16'b1111111110101011   ;
13'd1343:weight<=16'b0000000010010111   ;
13'd1344:weight<=16'b1111111110100111   ;
13'd1345:weight<=16'b1111111110011010   ;
13'd1346:weight<=16'b1111111111111000   ;
13'd1347:weight<=16'b0000000001011000   ;
13'd1348:weight<=16'b1111111111111010   ;
13'd1349:weight<=16'b0000000000010010   ;
13'd1350:weight<=16'b1111111100101011   ;
13'd1351:weight<=16'b0000010000011010   ;
13'd1352:weight<=16'b1111111110110010   ;
13'd1353:weight<=16'b1111111010110011   ;
13'd1354:weight<=16'b1111111100000000   ;
13'd1355:weight<=16'b0000000011101110   ;
13'd1356:weight<=16'b1111111101100001   ;
13'd1357:weight<=16'b1111111100110110   ;
13'd1358:weight<=16'b0000000001111101   ;
13'd1359:weight<=16'b0000000001001110   ;
13'd1360:weight<=16'b1111111111010000   ;
13'd1361:weight<=16'b0000000000000101   ;
13'd1362:weight<=16'b1111111110010110   ;
13'd1363:weight<=16'b0000000001000010   ;
13'd1364:weight<=16'b1111111111111011   ;
13'd1365:weight<=16'b0000000000011110   ;
13'd1366:weight<=16'b0000000011101000   ;
13'd1367:weight<=16'b0000000010110001   ;
13'd1368:weight<=16'b1111111110111000   ;
13'd1369:weight<=16'b1111111101001110   ;
13'd1370:weight<=16'b0000000001001011   ;
13'd1371:weight<=16'b0000000000000111   ;
13'd1372:weight<=16'b1111111111101110   ;
13'd1373:weight<=16'b1111111111111111   ;
13'd1374:weight<=16'b1111111111011000   ;
13'd1375:weight<=16'b1111111111111111   ;
13'd1376:weight<=16'b1111111111001110   ;
13'd1377:weight<=16'b0000000000111010   ;
13'd1378:weight<=16'b0000000001100000   ;
13'd1379:weight<=16'b1111111110110000   ;
13'd1380:weight<=16'b1111111110111011   ;
13'd1381:weight<=16'b1111111111010011   ;
13'd1382:weight<=16'b0000000000011010   ;
13'd1383:weight<=16'b1111111111011001   ;
13'd1384:weight<=16'b1111111100110011   ;
13'd1385:weight<=16'b1111111111011101   ;
13'd1386:weight<=16'b0000000100010011   ;
13'd1387:weight<=16'b0000000001111110   ;
13'd1388:weight<=16'b1111111111000100   ;
13'd1389:weight<=16'b0000000001001010   ;
13'd1390:weight<=16'b0000000011100111   ;
13'd1391:weight<=16'b1111111101111010   ;
13'd1392:weight<=16'b1111111110101011   ;
13'd1393:weight<=16'b0000000010010111   ;
13'd1394:weight<=16'b1111111110100111   ;
13'd1395:weight<=16'b1111111110011010   ;
13'd1396:weight<=16'b1111111111111000   ;
13'd1397:weight<=16'b0000000001011000   ;
13'd1398:weight<=16'b1111111111111010   ;
13'd1399:weight<=16'b0000000000010010   ;
13'd1400:weight<=16'b1111111110010100   ;
13'd1401:weight<=16'b1111111111001011   ;
13'd1402:weight<=16'b1111111111001001   ;
13'd1403:weight<=16'b0000000010000110   ;
13'd1404:weight<=16'b0000000100100101   ;
13'd1405:weight<=16'b0000000101010110   ;
13'd1406:weight<=16'b1111111111110011   ;
13'd1407:weight<=16'b1111111000101100   ;
13'd1408:weight<=16'b1111111000111001   ;
13'd1409:weight<=16'b0000000110100100   ;
13'd1410:weight<=16'b1111111111010000   ;
13'd1411:weight<=16'b0000000000000101   ;
13'd1412:weight<=16'b1111111110010110   ;
13'd1413:weight<=16'b0000000001000010   ;
13'd1414:weight<=16'b1111111111111011   ;
13'd1415:weight<=16'b0000000000011110   ;
13'd1416:weight<=16'b0000000011101000   ;
13'd1417:weight<=16'b0000000010110001   ;
13'd1418:weight<=16'b1111111110111000   ;
13'd1419:weight<=16'b1111111101001110   ;
13'd1420:weight<=16'b1111111111001000   ;
13'd1421:weight<=16'b0000000000010100   ;
13'd1422:weight<=16'b0000000000111110   ;
13'd1423:weight<=16'b0000000001001101   ;
13'd1424:weight<=16'b0000000001000011   ;
13'd1425:weight<=16'b1111111111101011   ;
13'd1426:weight<=16'b1111111101101011   ;
13'd1427:weight<=16'b1111111111001101   ;
13'd1428:weight<=16'b1111111111100100   ;
13'd1429:weight<=16'b0000000001010100   ;
13'd1430:weight<=16'b1111111110111011   ;
13'd1431:weight<=16'b1111111111010011   ;
13'd1432:weight<=16'b0000000000011010   ;
13'd1433:weight<=16'b1111111111011001   ;
13'd1434:weight<=16'b1111111100110011   ;
13'd1435:weight<=16'b1111111111011101   ;
13'd1436:weight<=16'b0000000100010011   ;
13'd1437:weight<=16'b0000000001111110   ;
13'd1438:weight<=16'b1111111111000100   ;
13'd1439:weight<=16'b0000000001001010   ;
13'd1440:weight<=16'b1111111110100100   ;
13'd1441:weight<=16'b0000000001110010   ;
13'd1442:weight<=16'b0000000010011011   ;
13'd1443:weight<=16'b0000000000100110   ;
13'd1444:weight<=16'b0000000000001110   ;
13'd1445:weight<=16'b1111111111011000   ;
13'd1446:weight<=16'b1111111111010011   ;
13'd1447:weight<=16'b1111111110001011   ;
13'd1448:weight<=16'b1111111111100001   ;
13'd1449:weight<=16'b0000000000110111   ;
13'd1450:weight<=16'b1111111110010100   ;
13'd1451:weight<=16'b1111111111001011   ;
13'd1452:weight<=16'b1111111111001001   ;
13'd1453:weight<=16'b0000000010000110   ;
13'd1454:weight<=16'b0000000100100101   ;
13'd1455:weight<=16'b0000000101010110   ;
13'd1456:weight<=16'b1111111111110011   ;
13'd1457:weight<=16'b1111111000101100   ;
13'd1458:weight<=16'b1111111000111001   ;
13'd1459:weight<=16'b0000000110100100   ;
13'd1460:weight<=16'b1111111111111001   ;
13'd1461:weight<=16'b0000000000110111   ;
13'd1462:weight<=16'b1111111111110000   ;
13'd1463:weight<=16'b0000000000011111   ;
13'd1464:weight<=16'b1111111111101101   ;
13'd1465:weight<=16'b0000000001000000   ;
13'd1466:weight<=16'b0000000001010000   ;
13'd1467:weight<=16'b1111111110110111   ;
13'd1468:weight<=16'b0000000000110010   ;
13'd1469:weight<=16'b1111111111011010   ;
13'd1470:weight<=16'b1111111111001000   ;
13'd1471:weight<=16'b0000000000010100   ;
13'd1472:weight<=16'b0000000000111110   ;
13'd1473:weight<=16'b0000000001001101   ;
13'd1474:weight<=16'b0000000001000011   ;
13'd1475:weight<=16'b1111111111101011   ;
13'd1476:weight<=16'b1111111101101011   ;
13'd1477:weight<=16'b1111111111001101   ;
13'd1478:weight<=16'b1111111111100100   ;
13'd1479:weight<=16'b0000000001010100   ;
13'd1480:weight<=16'b0000000001110001   ;
13'd1481:weight<=16'b0000000000100011   ;
13'd1482:weight<=16'b1111111110111010   ;
13'd1483:weight<=16'b1111111110101100   ;
13'd1484:weight<=16'b1111111111110100   ;
13'd1485:weight<=16'b1111111110010011   ;
13'd1486:weight<=16'b1111111110110100   ;
13'd1487:weight<=16'b1111111110101010   ;
13'd1488:weight<=16'b0000000001101011   ;
13'd1489:weight<=16'b0000000010101001   ;
13'd1490:weight<=16'b1111111110100100   ;
13'd1491:weight<=16'b0000000001110010   ;
13'd1492:weight<=16'b0000000010011011   ;
13'd1493:weight<=16'b0000000000100110   ;
13'd1494:weight<=16'b0000000000001110   ;
13'd1495:weight<=16'b1111111111011000   ;
13'd1496:weight<=16'b1111111111010011   ;
13'd1497:weight<=16'b1111111110001011   ;
13'd1498:weight<=16'b1111111111100001   ;
13'd1499:weight<=16'b0000000000110111   ;
13'd1500:weight<=16'b0000000110101000   ;
13'd1501:weight<=16'b1111111110110111   ;
13'd1502:weight<=16'b0000000010011000   ;
13'd1503:weight<=16'b1111111000100011   ;
13'd1504:weight<=16'b1111111101100111   ;
13'd1505:weight<=16'b1111111111011000   ;
13'd1506:weight<=16'b1111111101000101   ;
13'd1507:weight<=16'b0000000001101011   ;
13'd1508:weight<=16'b0000000000000110   ;
13'd1509:weight<=16'b0000000100110100   ;
13'd1510:weight<=16'b1111111111111001   ;
13'd1511:weight<=16'b0000000000110111   ;
13'd1512:weight<=16'b1111111111110000   ;
13'd1513:weight<=16'b0000000000011111   ;
13'd1514:weight<=16'b1111111111101101   ;
13'd1515:weight<=16'b0000000001000000   ;
13'd1516:weight<=16'b0000000001010000   ;
13'd1517:weight<=16'b1111111110110111   ;
13'd1518:weight<=16'b0000000000110010   ;
13'd1519:weight<=16'b1111111111011010   ;
13'd1520:weight<=16'b0000000000001100   ;
13'd1521:weight<=16'b0000000000011001   ;
13'd1522:weight<=16'b1111111100010111   ;
13'd1523:weight<=16'b0000000001010001   ;
13'd1524:weight<=16'b0000000000111000   ;
13'd1525:weight<=16'b0000000000000100   ;
13'd1526:weight<=16'b1111111111100011   ;
13'd1527:weight<=16'b1111111111010000   ;
13'd1528:weight<=16'b0000000010000101   ;
13'd1529:weight<=16'b0000000000111001   ;
13'd1530:weight<=16'b0000000001110001   ;
13'd1531:weight<=16'b0000000000100011   ;
13'd1532:weight<=16'b1111111110111010   ;
13'd1533:weight<=16'b1111111110101100   ;
13'd1534:weight<=16'b1111111111110100   ;
13'd1535:weight<=16'b1111111110010011   ;
13'd1536:weight<=16'b1111111110110100   ;
13'd1537:weight<=16'b1111111110101010   ;
13'd1538:weight<=16'b0000000001101011   ;
13'd1539:weight<=16'b0000000010101001   ;
13'd1540:weight<=16'b1111111111111110   ;
13'd1541:weight<=16'b1111111111110111   ;
13'd1542:weight<=16'b1111111110101101   ;
13'd1543:weight<=16'b0000000000001111   ;
13'd1544:weight<=16'b1111111111111101   ;
13'd1545:weight<=16'b1111111111000111   ;
13'd1546:weight<=16'b0000000010001000   ;
13'd1547:weight<=16'b1111111111100011   ;
13'd1548:weight<=16'b0000000000101111   ;
13'd1549:weight<=16'b1111111111111101   ;
13'd1550:weight<=16'b0000000110101000   ;
13'd1551:weight<=16'b1111111110110111   ;
13'd1552:weight<=16'b0000000010011000   ;
13'd1553:weight<=16'b1111111000100011   ;
13'd1554:weight<=16'b1111111101100111   ;
13'd1555:weight<=16'b1111111111011000   ;
13'd1556:weight<=16'b1111111101000101   ;
13'd1557:weight<=16'b0000000001101011   ;
13'd1558:weight<=16'b0000000000000110   ;
13'd1559:weight<=16'b0000000100110100   ;
13'd1560:weight<=16'b1111111111100001   ;
13'd1561:weight<=16'b1111111111010110   ;
13'd1562:weight<=16'b0000000000101000   ;
13'd1563:weight<=16'b0000000010011010   ;
13'd1564:weight<=16'b0000000000110101   ;
13'd1565:weight<=16'b0000000000011000   ;
13'd1566:weight<=16'b0000000000100100   ;
13'd1567:weight<=16'b1111111110001011   ;
13'd1568:weight<=16'b1111111111100001   ;
13'd1569:weight<=16'b1111111111110001   ;
13'd1570:weight<=16'b0000000000001100   ;
13'd1571:weight<=16'b0000000000011001   ;
13'd1572:weight<=16'b1111111100010111   ;
13'd1573:weight<=16'b0000000001010001   ;
13'd1574:weight<=16'b0000000000111000   ;
13'd1575:weight<=16'b0000000000000100   ;
13'd1576:weight<=16'b1111111111100011   ;
13'd1577:weight<=16'b1111111111010000   ;
13'd1578:weight<=16'b0000000010000101   ;
13'd1579:weight<=16'b0000000000111001   ;
13'd1580:weight<=16'b0000000000000101   ;
13'd1581:weight<=16'b0000000000001110   ;
13'd1582:weight<=16'b1111111101111010   ;
13'd1583:weight<=16'b1111111110001111   ;
13'd1584:weight<=16'b1111111111010000   ;
13'd1585:weight<=16'b1111111111000100   ;
13'd1586:weight<=16'b0000000010011001   ;
13'd1587:weight<=16'b0000000000101000   ;
13'd1588:weight<=16'b0000000000011110   ;
13'd1589:weight<=16'b0000000001101110   ;
13'd1590:weight<=16'b1111111111111110   ;
13'd1591:weight<=16'b1111111111110111   ;
13'd1592:weight<=16'b1111111110101101   ;
13'd1593:weight<=16'b0000000000001111   ;
13'd1594:weight<=16'b1111111111111101   ;
13'd1595:weight<=16'b1111111111000111   ;
13'd1596:weight<=16'b0000000010001000   ;
13'd1597:weight<=16'b1111111111100011   ;
13'd1598:weight<=16'b0000000000101111   ;
13'd1599:weight<=16'b1111111111111101   ;
13'd1600:weight<=16'b0000000000101001   ;
13'd1601:weight<=16'b0000000000111110   ;
13'd1602:weight<=16'b0000000000011111   ;
13'd1603:weight<=16'b1111111111010100   ;
13'd1604:weight<=16'b1111111110001000   ;
13'd1605:weight<=16'b1111111111111111   ;
13'd1606:weight<=16'b0000000001001101   ;
13'd1607:weight<=16'b1111111101111001   ;
13'd1608:weight<=16'b1111111111100111   ;
13'd1609:weight<=16'b0000000010001001   ;
13'd1610:weight<=16'b1111111111100001   ;
13'd1611:weight<=16'b1111111111010110   ;
13'd1612:weight<=16'b0000000000101000   ;
13'd1613:weight<=16'b0000000010011010   ;
13'd1614:weight<=16'b0000000000110101   ;
13'd1615:weight<=16'b0000000000011000   ;
13'd1616:weight<=16'b0000000000100100   ;
13'd1617:weight<=16'b1111111110001011   ;
13'd1618:weight<=16'b1111111111100001   ;
13'd1619:weight<=16'b1111111111110001   ;
13'd1620:weight<=16'b0000000011000101   ;
13'd1621:weight<=16'b0000001000110111   ;
13'd1622:weight<=16'b1111111011100010   ;
13'd1623:weight<=16'b0000000101001010   ;
13'd1624:weight<=16'b1111111000011001   ;
13'd1625:weight<=16'b0000000001111011   ;
13'd1626:weight<=16'b1111111111011000   ;
13'd1627:weight<=16'b0000000000000011   ;
13'd1628:weight<=16'b1111111111100001   ;
13'd1629:weight<=16'b1111111100000111   ;
13'd1630:weight<=16'b0000000000000101   ;
13'd1631:weight<=16'b0000000000001110   ;
13'd1632:weight<=16'b1111111101111010   ;
13'd1633:weight<=16'b1111111110001111   ;
13'd1634:weight<=16'b1111111111010000   ;
13'd1635:weight<=16'b1111111111000100   ;
13'd1636:weight<=16'b0000000010011001   ;
13'd1637:weight<=16'b0000000000101000   ;
13'd1638:weight<=16'b0000000000011110   ;
13'd1639:weight<=16'b0000000001101110   ;
13'd1640:weight<=16'b1111111110110110   ;
13'd1641:weight<=16'b1111111101100011   ;
13'd1642:weight<=16'b0000000000110001   ;
13'd1643:weight<=16'b1111111111011000   ;
13'd1644:weight<=16'b0000000010011100   ;
13'd1645:weight<=16'b0000000010000011   ;
13'd1646:weight<=16'b1111111110101100   ;
13'd1647:weight<=16'b1111111110111110   ;
13'd1648:weight<=16'b0000000001100001   ;
13'd1649:weight<=16'b1111111111110110   ;
13'd1650:weight<=16'b0000000000101001   ;
13'd1651:weight<=16'b0000000000111110   ;
13'd1652:weight<=16'b0000000000011111   ;
13'd1653:weight<=16'b1111111111010100   ;
13'd1654:weight<=16'b1111111110001000   ;
13'd1655:weight<=16'b1111111111111111   ;
13'd1656:weight<=16'b0000000001001101   ;
13'd1657:weight<=16'b1111111101111001   ;
13'd1658:weight<=16'b1111111111100111   ;
13'd1659:weight<=16'b0000000010001001   ;
13'd1660:weight<=16'b1111111110111011   ;
13'd1661:weight<=16'b0000000000010010   ;
13'd1662:weight<=16'b1111111110111000   ;
13'd1663:weight<=16'b1111111111111011   ;
13'd1664:weight<=16'b0000000000100100   ;
13'd1665:weight<=16'b1111111111001011   ;
13'd1666:weight<=16'b0000000100011000   ;
13'd1667:weight<=16'b1111111111111111   ;
13'd1668:weight<=16'b1111111111000000   ;
13'd1669:weight<=16'b1111111111001111   ;
13'd1670:weight<=16'b0000000011000101   ;
13'd1671:weight<=16'b0000001000110111   ;
13'd1672:weight<=16'b1111111011100010   ;
13'd1673:weight<=16'b0000000101001010   ;
13'd1674:weight<=16'b1111111000011001   ;
13'd1675:weight<=16'b0000000001111011   ;
13'd1676:weight<=16'b1111111111011000   ;
13'd1677:weight<=16'b0000000000000011   ;
13'd1678:weight<=16'b1111111111100001   ;
13'd1679:weight<=16'b1111111100000111   ;
13'd1680:weight<=16'b0000000010010110   ;
13'd1681:weight<=16'b0000000000001111   ;
13'd1682:weight<=16'b1111111010111010   ;
13'd1683:weight<=16'b0000000011100010   ;
13'd1684:weight<=16'b0000000000110101   ;
13'd1685:weight<=16'b0000001000010110   ;
13'd1686:weight<=16'b1111111101111101   ;
13'd1687:weight<=16'b1111111110000010   ;
13'd1688:weight<=16'b1111111110111111   ;
13'd1689:weight<=16'b1111111100011011   ;
13'd1690:weight<=16'b1111111110110110   ;
13'd1691:weight<=16'b1111111101100011   ;
13'd1692:weight<=16'b0000000000110001   ;
13'd1693:weight<=16'b1111111111011000   ;
13'd1694:weight<=16'b0000000010011100   ;
13'd1695:weight<=16'b0000000010000011   ;
13'd1696:weight<=16'b1111111110101100   ;
13'd1697:weight<=16'b1111111110111110   ;
13'd1698:weight<=16'b0000000001100001   ;
13'd1699:weight<=16'b1111111111110110   ;
13'd1700:weight<=16'b0000000000001110   ;
13'd1701:weight<=16'b0000000000111000   ;
13'd1702:weight<=16'b0000000001111111   ;
13'd1703:weight<=16'b0000000010010100   ;
13'd1704:weight<=16'b1111111111010111   ;
13'd1705:weight<=16'b1111111110010101   ;
13'd1706:weight<=16'b0000000000001101   ;
13'd1707:weight<=16'b0000000001000000   ;
13'd1708:weight<=16'b1111111111111110   ;
13'd1709:weight<=16'b1111111101100111   ;
13'd1710:weight<=16'b1111111110111011   ;
13'd1711:weight<=16'b0000000000010010   ;
13'd1712:weight<=16'b1111111110111000   ;
13'd1713:weight<=16'b1111111111111011   ;
13'd1714:weight<=16'b0000000000100100   ;
13'd1715:weight<=16'b1111111111001011   ;
13'd1716:weight<=16'b0000000100011000   ;
13'd1717:weight<=16'b1111111111111111   ;
13'd1718:weight<=16'b1111111111000000   ;
13'd1719:weight<=16'b1111111111001111   ;
13'd1720:weight<=16'b0000000001001111   ;
13'd1721:weight<=16'b0000000001010011   ;
13'd1722:weight<=16'b0000000010110000   ;
13'd1723:weight<=16'b1111111110110110   ;
13'd1724:weight<=16'b0000000001000010   ;
13'd1725:weight<=16'b0000000001011000   ;
13'd1726:weight<=16'b1111111011001111   ;
13'd1727:weight<=16'b0000000001010001   ;
13'd1728:weight<=16'b1111111111101110   ;
13'd1729:weight<=16'b1111111110101000   ;
13'd1730:weight<=16'b0000000010010110   ;
13'd1731:weight<=16'b0000000000001111   ;
13'd1732:weight<=16'b1111111010111010   ;
13'd1733:weight<=16'b0000000011100010   ;
13'd1734:weight<=16'b0000000000110101   ;
13'd1735:weight<=16'b0000001000010110   ;
13'd1736:weight<=16'b1111111101111101   ;
13'd1737:weight<=16'b1111111110000010   ;
13'd1738:weight<=16'b1111111110111111   ;
13'd1739:weight<=16'b1111111100011011   ;
13'd1740:weight<=16'b0000000000001010   ;
13'd1741:weight<=16'b0000000001110011   ;
13'd1742:weight<=16'b1111111110001101   ;
13'd1743:weight<=16'b0000000000001110   ;
13'd1744:weight<=16'b1111111110110011   ;
13'd1745:weight<=16'b0000000000100001   ;
13'd1746:weight<=16'b1111111110011011   ;
13'd1747:weight<=16'b0000000000010111   ;
13'd1748:weight<=16'b0000000000101111   ;
13'd1749:weight<=16'b0000000001000000   ;
13'd1750:weight<=16'b0000000000001110   ;
13'd1751:weight<=16'b0000000000111000   ;
13'd1752:weight<=16'b0000000001111111   ;
13'd1753:weight<=16'b0000000010010100   ;
13'd1754:weight<=16'b1111111111010111   ;
13'd1755:weight<=16'b1111111110010101   ;
13'd1756:weight<=16'b0000000000001101   ;
13'd1757:weight<=16'b0000000001000000   ;
13'd1758:weight<=16'b1111111111111110   ;
13'd1759:weight<=16'b1111111101100111   ;
13'd1760:weight<=16'b1111111110011110   ;
13'd1761:weight<=16'b1111111101110110   ;
13'd1762:weight<=16'b1111111101000011   ;
13'd1763:weight<=16'b0000000100011010   ;
13'd1764:weight<=16'b1111111110101111   ;
13'd1765:weight<=16'b0000000001001100   ;
13'd1766:weight<=16'b0000000000111001   ;
13'd1767:weight<=16'b0000000001110010   ;
13'd1768:weight<=16'b0000000000001100   ;
13'd1769:weight<=16'b0000000000010110   ;
13'd1770:weight<=16'b0000000001001111   ;
13'd1771:weight<=16'b0000000001010011   ;
13'd1772:weight<=16'b0000000010110000   ;
13'd1773:weight<=16'b1111111110110110   ;
13'd1774:weight<=16'b0000000001000010   ;
13'd1775:weight<=16'b0000000001011000   ;
13'd1776:weight<=16'b1111111011001111   ;
13'd1777:weight<=16'b0000000001010001   ;
13'd1778:weight<=16'b1111111111101110   ;
13'd1779:weight<=16'b1111111110101000   ;
13'd1780:weight<=16'b1111111110110100   ;
13'd1781:weight<=16'b0000000101011110   ;
13'd1782:weight<=16'b1111111111010000   ;
13'd1783:weight<=16'b1111111111111101   ;
13'd1784:weight<=16'b0000000011101001   ;
13'd1785:weight<=16'b1111111111001011   ;
13'd1786:weight<=16'b1111111110110011   ;
13'd1787:weight<=16'b1111111101101100   ;
13'd1788:weight<=16'b1111111111111111   ;
13'd1789:weight<=16'b1111111111001010   ;
13'd1790:weight<=16'b0000000000001010   ;
13'd1791:weight<=16'b0000000001110011   ;
13'd1792:weight<=16'b1111111110001101   ;
13'd1793:weight<=16'b0000000000001110   ;
13'd1794:weight<=16'b1111111110110011   ;
13'd1795:weight<=16'b0000000000100001   ;
13'd1796:weight<=16'b1111111110011011   ;
13'd1797:weight<=16'b0000000000010111   ;
13'd1798:weight<=16'b0000000000101111   ;
13'd1799:weight<=16'b0000000001000000   ;
13'd1800:weight<=16'b0000000000011111   ;
13'd1801:weight<=16'b1111111111000000   ;
13'd1802:weight<=16'b0000000011110001   ;
13'd1803:weight<=16'b1111111110011110   ;
13'd1804:weight<=16'b1111111110011001   ;
13'd1805:weight<=16'b0000000010101000   ;
13'd1806:weight<=16'b1111111111101001   ;
13'd1807:weight<=16'b1111111111111110   ;
13'd1808:weight<=16'b1111111111000111   ;
13'd1809:weight<=16'b1111111111101110   ;
13'd1810:weight<=16'b1111111110011110   ;
13'd1811:weight<=16'b1111111101110110   ;
13'd1812:weight<=16'b1111111101000011   ;
13'd1813:weight<=16'b0000000100011010   ;
13'd1814:weight<=16'b1111111110101111   ;
13'd1815:weight<=16'b0000000001001100   ;
13'd1816:weight<=16'b0000000000111001   ;
13'd1817:weight<=16'b0000000001110010   ;
13'd1818:weight<=16'b0000000000001100   ;
13'd1819:weight<=16'b0000000000010110   ;
13'd1820:weight<=16'b0000000001011111   ;
13'd1821:weight<=16'b1111111110110011   ;
13'd1822:weight<=16'b1111111111100111   ;
13'd1823:weight<=16'b1111111110010010   ;
13'd1824:weight<=16'b1111111110111101   ;
13'd1825:weight<=16'b1111111110001001   ;
13'd1826:weight<=16'b0000000010100001   ;
13'd1827:weight<=16'b0000000100110001   ;
13'd1828:weight<=16'b1111111111101010   ;
13'd1829:weight<=16'b1111111111010000   ;
13'd1830:weight<=16'b1111111110110100   ;
13'd1831:weight<=16'b0000000101011110   ;
13'd1832:weight<=16'b1111111111010000   ;
13'd1833:weight<=16'b1111111111111101   ;
13'd1834:weight<=16'b0000000011101001   ;
13'd1835:weight<=16'b1111111111001011   ;
13'd1836:weight<=16'b1111111110110011   ;
13'd1837:weight<=16'b1111111101101100   ;
13'd1838:weight<=16'b1111111111111111   ;
13'd1839:weight<=16'b1111111111001010   ;
13'd1840:weight<=16'b1111111111111000   ;
13'd1841:weight<=16'b0000000001101110   ;
13'd1842:weight<=16'b0000000010101100   ;
13'd1843:weight<=16'b0000000000100101   ;
13'd1844:weight<=16'b1111111110110001   ;
13'd1845:weight<=16'b1111111111110110   ;
13'd1846:weight<=16'b0000000011010000   ;
13'd1847:weight<=16'b1111111111100101   ;
13'd1848:weight<=16'b1111111000101111   ;
13'd1849:weight<=16'b0000000010101001   ;
13'd1850:weight<=16'b0000000000011111   ;
13'd1851:weight<=16'b1111111111000000   ;
13'd1852:weight<=16'b0000000011110001   ;
13'd1853:weight<=16'b1111111110011110   ;
13'd1854:weight<=16'b1111111110011001   ;
13'd1855:weight<=16'b0000000010101000   ;
13'd1856:weight<=16'b1111111111101001   ;
13'd1857:weight<=16'b1111111111111110   ;
13'd1858:weight<=16'b1111111111000111   ;
13'd1859:weight<=16'b1111111111101110   ;
13'd1860:weight<=16'b1111111111000101   ;
13'd1861:weight<=16'b1111111111111101   ;
13'd1862:weight<=16'b1111111110100110   ;
13'd1863:weight<=16'b0000000011100000   ;
13'd1864:weight<=16'b1111111111101111   ;
13'd1865:weight<=16'b0000000000101000   ;
13'd1866:weight<=16'b1111111111110101   ;
13'd1867:weight<=16'b1111111111110100   ;
13'd1868:weight<=16'b1111111111110001   ;
13'd1869:weight<=16'b1111111111011111  ;
13'd1870:weight<=16'b0000000001011111   ;
13'd1871:weight<=16'b1111111110110011   ;
13'd1872:weight<=16'b1111111111100111   ;
13'd1873:weight<=16'b1111111110010010   ;
13'd1874:weight<=16'b1111111110111101   ;
13'd1875:weight<=16'b1111111110001001   ;
13'd1876:weight<=16'b0000000010100001   ;
13'd1877:weight<=16'b0000000100110001   ;
13'd1878:weight<=16'b1111111111101010   ;
13'd1879:weight<=16'b1111111111010000   ;
13'd1880:weight<=16'b1111111111010111   ;
13'd1881:weight<=16'b1111111111101111   ;
13'd1882:weight<=16'b0000000000010100   ;
13'd1883:weight<=16'b1111111111100111   ;
13'd1884:weight<=16'b1111111111011011   ;
13'd1885:weight<=16'b1111111110101110   ;
13'd1886:weight<=16'b0000000001001011   ;
13'd1887:weight<=16'b0000000001110011   ;
13'd1888:weight<=16'b0000000000010000   ;
13'd1889:weight<=16'b1111111111100111   ;
13'd1890:weight<=16'b1111111111111000   ;
13'd1891:weight<=16'b0000000001101110   ;
13'd1892:weight<=16'b0000000010101100   ;
13'd1893:weight<=16'b0000000000100101   ;
13'd1894:weight<=16'b1111111110110001   ;
13'd1895:weight<=16'b1111111111110110   ;
13'd1896:weight<=16'b0000000011010000   ;
13'd1897:weight<=16'b1111111111100101   ;
13'd1898:weight<=16'b1111111000101111   ;
13'd1899:weight<=16'b0000000010101001   ;
13'd1900:weight<=16'b0000000000001110   ;
13'd1901:weight<=16'b1111111110000001   ;
13'd1902:weight<=16'b1111111111110110   ;
13'd1903:weight<=16'b1111111101110111   ;
13'd1904:weight<=16'b0000000001011000   ;
13'd1905:weight<=16'b0000000001011011   ;
13'd1906:weight<=16'b1111111111101101   ;
13'd1907:weight<=16'b0000000001001111   ;
13'd1908:weight<=16'b0000000001110111   ;
13'd1909:weight<=16'b1111111110111110   ;
13'd1910:weight<=16'b1111111111000101   ;
13'd1911:weight<=16'b1111111111111101   ;
13'd1912:weight<=16'b1111111110100110   ;
13'd1913:weight<=16'b0000000011100000   ;
13'd1914:weight<=16'b1111111111101111   ;
13'd1915:weight<=16'b0000000000101000   ;
13'd1916:weight<=16'b1111111111110101   ;
13'd1917:weight<=16'b1111111111110100   ;
13'd1918:weight<=16'b1111111111110001   ;
13'd1919:weight<=16'b1111111111011111   ;
13'd1920:weight<=16'b0000000000110001   ;
13'd1921:weight<=16'b1111111110011110   ;
13'd1922:weight<=16'b0000000000000011   ;
13'd1923:weight<=16'b0000000100110100   ;
13'd1924:weight<=16'b1111111101010101   ;
13'd1925:weight<=16'b1111111100011110   ;
13'd1926:weight<=16'b0000000000010000   ;
13'd1927:weight<=16'b0000000010010010   ;
13'd1928:weight<=16'b0000000001000101   ;
13'd1929:weight<=16'b1111111111100001   ;
13'd1930:weight<=16'b1111111111010111   ;
13'd1931:weight<=16'b1111111111101111   ;
13'd1932:weight<=16'b0000000000010100   ;
13'd1933:weight<=16'b1111111111100111   ;
13'd1934:weight<=16'b1111111111011011   ;
13'd1935:weight<=16'b1111111110101110   ;
13'd1936:weight<=16'b0000000001001011   ;
13'd1937:weight<=16'b0000000001110011   ;
13'd1938:weight<=16'b0000000000010000   ;
13'd1939:weight<=16'b1111111111100111   ;
13'd1940:weight<=16'b1111111110101001   ;
13'd1941:weight<=16'b0000000100100110   ;
13'd1942:weight<=16'b0000000001001000   ;
13'd1943:weight<=16'b1111111111100010   ;
13'd1944:weight<=16'b0000000000101010   ;
13'd1945:weight<=16'b1111111111110101   ;
13'd1946:weight<=16'b0000000000000010   ;
13'd1947:weight<=16'b1111111101110000   ;
13'd1948:weight<=16'b1111111101100110   ;
13'd1949:weight<=16'b0000000000010101   ;
13'd1950:weight<=16'b0000000000001110   ;
13'd1951:weight<=16'b1111111110000001   ;
13'd1952:weight<=16'b1111111111110110   ;
13'd1953:weight<=16'b1111111101110111   ;
13'd1954:weight<=16'b0000000001011000   ;
13'd1955:weight<=16'b0000000001011011   ;
13'd1956:weight<=16'b1111111111101101   ;
13'd1957:weight<=16'b0000000001001111   ;
13'd1958:weight<=16'b0000000001110111   ;
13'd1959:weight<=16'b1111111110111110   ;
13'd1960:weight<=16'b0000000000000111   ;
13'd1961:weight<=16'b0000000001010000   ;
13'd1962:weight<=16'b0000000001010001   ;
13'd1963:weight<=16'b0000000001111101   ;
13'd1964:weight<=16'b1111111111111110   ;
13'd1965:weight<=16'b1111111101011110   ;
13'd1966:weight<=16'b1111111111100010   ;
13'd1967:weight<=16'b0000000000010101   ;
13'd1968:weight<=16'b0000000000000010   ;
13'd1969:weight<=16'b1111111111001111   ;
13'd1970:weight<=16'b0000000000110001   ;
13'd1971:weight<=16'b1111111110011110   ;
13'd1972:weight<=16'b0000000000000011   ;
13'd1973:weight<=16'b0000000100110100   ;
13'd1974:weight<=16'b1111111101010101   ;
13'd1975:weight<=16'b1111111100011110   ;
13'd1976:weight<=16'b0000000000010000   ;
13'd1977:weight<=16'b0000000010010010   ;
13'd1978:weight<=16'b0000000001000101   ;
13'd1979:weight<=16'b1111111111100001   ;
13'd1980:weight<=16'b0000000000000010   ;
13'd1981:weight<=16'b0000000000001101   ;
13'd1982:weight<=16'b0000000010000000   ;
13'd1983:weight<=16'b1111111101011110   ;
13'd1984:weight<=16'b1111111111111100   ;
13'd1985:weight<=16'b0000000001110111   ;
13'd1986:weight<=16'b0000000010000000   ;
13'd1987:weight<=16'b0000000000010100   ;
13'd1988:weight<=16'b1111111110000001   ;
13'd1989:weight<=16'b1111111110110110   ;
13'd1990:weight<=16'b1111111110101001   ;
13'd1991:weight<=16'b0000000100100110   ;
13'd1992:weight<=16'b0000000001001000   ;
13'd1993:weight<=16'b1111111111100010   ;
13'd1994:weight<=16'b0000000000101010   ;
13'd1995:weight<=16'b1111111111110101   ;
13'd1996:weight<=16'b0000000000000010   ;
13'd1997:weight<=16'b1111111101110000   ;
13'd1998:weight<=16'b1111111101100110   ;
13'd1999:weight<=16'b0000000000010101   ;
13'd2000:weight<=16'b1111111111001111   ;
13'd2001:weight<=16'b0000000001010101   ;
13'd2002:weight<=16'b1111111111000000   ;
13'd2003:weight<=16'b1111111111011000   ;
13'd2004:weight<=16'b0000000000110101   ;
13'd2005:weight<=16'b1111111110111110   ;
13'd2006:weight<=16'b1111111111101100   ;
13'd2007:weight<=16'b1111111111011011   ;
13'd2008:weight<=16'b0000000000111010   ;
13'd2009:weight<=16'b0000000001110100   ;
13'd2010:weight<=16'b0000000000000111   ;
13'd2011:weight<=16'b0000000001010000   ;
13'd2012:weight<=16'b0000000001010001   ;
13'd2013:weight<=16'b0000000001111101   ;
13'd2014:weight<=16'b1111111111111110   ;
13'd2015:weight<=16'b1111111101011110  ;
13'd2016:weight<=16'b1111111111100010   ;
13'd2017:weight<=16'b0000000000010101   ;
13'd2018:weight<=16'b0000000000000010   ;
13'd2019:weight<=16'b1111111111001111   ;
13'd2020:weight<=16'b1111111011110010   ;
13'd2021:weight<=16'b1111111000010010   ;
13'd2022:weight<=16'b0000000011110001   ;
13'd2023:weight<=16'b1111111111100011   ;
13'd2024:weight<=16'b0000000011110110   ;
13'd2025:weight<=16'b1111111110000000   ;
13'd2026:weight<=16'b1111111111010001   ;
13'd2027:weight<=16'b0000000100100111   ;
13'd2028:weight<=16'b1111111101111101   ;
13'd2029:weight<=16'b0000000110101011   ;
13'd2030:weight<=16'b0000000000000010   ;
13'd2031:weight<=16'b0000000000001101   ;
13'd2032:weight<=16'b0000000010000000   ;
13'd2033:weight<=16'b1111111101011110   ;
13'd2034:weight<=16'b1111111111111100   ;
13'd2035:weight<=16'b0000000001110111   ;
13'd2036:weight<=16'b0000000010000000   ;
13'd2037:weight<=16'b0000000000010100   ;
13'd2038:weight<=16'b1111111110000001   ;
13'd2039:weight<=16'b1111111110110110   ;
13'd2040:weight<=16'b1111111111000110   ;
13'd2041:weight<=16'b1111111111100000   ;
13'd2042:weight<=16'b1111111110010010   ;
13'd2043:weight<=16'b0000000010011100   ;
13'd2044:weight<=16'b0000000001101000   ;
13'd2045:weight<=16'b1111111111010000   ;
13'd2046:weight<=16'b1111111111110111   ;
13'd2047:weight<=16'b0000000000100000   ;
13'd2048:weight<=16'b1111111111111001   ;
13'd2049:weight<=16'b1111111111011011   ;
13'd2050:weight<=16'b1111111111001111   ;
13'd2051:weight<=16'b0000000001010101   ;
13'd2052:weight<=16'b1111111111000000   ;
13'd2053:weight<=16'b1111111111011000   ;
13'd2054:weight<=16'b0000000000110101   ;
13'd2055:weight<=16'b1111111110111110   ;
13'd2056:weight<=16'b1111111111101100   ;
13'd2057:weight<=16'b1111111111011011   ;
13'd2058:weight<=16'b0000000000111010   ;
13'd2059:weight<=16'b0000000001110100   ;
13'd2060:weight<=16'b1111111111110010   ;
13'd2061:weight<=16'b1111111101111000   ;
13'd2062:weight<=16'b1111111110101011   ;
13'd2063:weight<=16'b0000000010100111   ;
13'd2064:weight<=16'b0000000001001111   ;
13'd2065:weight<=16'b0000000000101011   ;
13'd2066:weight<=16'b1111111111001110   ;
13'd2067:weight<=16'b0000000001010100   ;
13'd2068:weight<=16'b0000000001101000   ;
13'd2069:weight<=16'b1111111110101000   ;
13'd2070:weight<=16'b1111111011110010   ;
13'd2071:weight<=16'b1111111000010010   ;
13'd2072:weight<=16'b0000000011110001   ;
13'd2073:weight<=16'b1111111111100011   ;
13'd2074:weight<=16'b0000000011110110   ;
13'd2075:weight<=16'b1111111110000000   ;
13'd2076:weight<=16'b1111111111010001   ;
13'd2077:weight<=16'b0000000100100111   ;
13'd2078:weight<=16'b1111111101111101   ;
13'd2079:weight<=16'b0000000110101011   ;
13'd2080:weight<=16'b0000000001000000   ;
13'd2081:weight<=16'b1111111111101001   ;
13'd2082:weight<=16'b1111111100111100   ;
13'd2083:weight<=16'b1111111111010111   ;
13'd2084:weight<=16'b1111111100111101   ;
13'd2085:weight<=16'b0000000000010111   ;
13'd2086:weight<=16'b0000000000111001   ;
13'd2087:weight<=16'b0000000011010010   ;
13'd2088:weight<=16'b0000000010010010   ;
13'd2089:weight<=16'b0000000000001000   ;
13'd2090:weight<=16'b1111111111000110   ;
13'd2091:weight<=16'b1111111111100000   ;
13'd2092:weight<=16'b1111111110010010   ;
13'd2093:weight<=16'b0000000010011100   ;
13'd2094:weight<=16'b0000000001101000   ;
13'd2095:weight<=16'b1111111111010000   ;
13'd2096:weight<=16'b1111111111110111   ;
13'd2097:weight<=16'b0000000000100000   ;
13'd2098:weight<=16'b1111111111111001   ;
13'd2099:weight<=16'b1111111111011011   ;
13'd2100:weight<=16'b1111111110110101   ;
13'd2101:weight<=16'b1111111111111000   ;
13'd2102:weight<=16'b1111111110110000   ;
13'd2103:weight<=16'b0000000000111111   ;
13'd2104:weight<=16'b0000000000000101   ;
13'd2105:weight<=16'b0000000010001001   ;
13'd2106:weight<=16'b1111111110010001   ;
13'd2107:weight<=16'b0000000001111111   ;
13'd2108:weight<=16'b1111111111000110   ;
13'd2109:weight<=16'b0000000000010100   ;
13'd2110:weight<=16'b1111111111110010   ;
13'd2111:weight<=16'b1111111101111000   ;
13'd2112:weight<=16'b1111111110101011   ;
13'd2113:weight<=16'b0000000010100111   ;
13'd2114:weight<=16'b0000000001001111   ;
13'd2115:weight<=16'b0000000000101011   ;
13'd2116:weight<=16'b1111111111001110   ;
13'd2117:weight<=16'b0000000001010100   ;
13'd2118:weight<=16'b0000000001101000   ;
13'd2119:weight<=16'b1111111110101000   ;
13'd2120:weight<=16'b1111111111100000   ;
13'd2121:weight<=16'b0000001000101000   ;
13'd2122:weight<=16'b1111111101111010   ;
13'd2123:weight<=16'b0000000101011101   ;
13'd2124:weight<=16'b0000010101111000   ;
13'd2125:weight<=16'b0000010100000110   ;
13'd2126:weight<=16'b1111101011010011   ;
13'd2127:weight<=16'b1111101001101101   ;
13'd2128:weight<=16'b1111110111010000   ;
13'd2129:weight<=16'b0000000100001111   ;
13'd2130:weight<=16'b0000000001000000   ;
13'd2131:weight<=16'b1111111111101001   ;
13'd2132:weight<=16'b1111111100111100   ;
13'd2133:weight<=16'b1111111111010111   ;
13'd2134:weight<=16'b1111111100111101   ;
13'd2135:weight<=16'b0000000000010111   ;
13'd2136:weight<=16'b0000000000111001   ;
13'd2137:weight<=16'b0000000011010010   ;
13'd2138:weight<=16'b0000000010010010   ;
13'd2139:weight<=16'b0000000000001000   ;
13'd2140:weight<=16'b1111111111000100   ;
13'd2141:weight<=16'b1111111111100111   ;
13'd2142:weight<=16'b1111111111100011   ;
13'd2143:weight<=16'b1111111110100101   ;
13'd2144:weight<=16'b0000000000100010   ;
13'd2145:weight<=16'b1111111111101111   ;
13'd2146:weight<=16'b0000000001000011   ;
13'd2147:weight<=16'b0000000001010000   ;
13'd2148:weight<=16'b1111111111100111   ;
13'd2149:weight<=16'b0000000001100011   ;
13'd2150:weight<=16'b1111111110110101   ;
13'd2151:weight<=16'b1111111111111000   ;
13'd2152:weight<=16'b1111111110110000   ;
13'd2153:weight<=16'b0000000000111111   ;
13'd2154:weight<=16'b0000000000000101   ;
13'd2155:weight<=16'b0000000010001001   ;
13'd2156:weight<=16'b1111111110010001   ;
13'd2157:weight<=16'b0000000001111111   ;
13'd2158:weight<=16'b1111111111000110   ;
13'd2159:weight<=16'b0000000000010100   ;
13'd2160:weight<=16'b1111111101100100   ;
13'd2161:weight<=16'b1111111110001111   ;
13'd2162:weight<=16'b1111111111000011   ;
13'd2163:weight<=16'b0000000000110110   ;
13'd2164:weight<=16'b1111111111100010   ;
13'd2165:weight<=16'b0000000000111011   ;
13'd2166:weight<=16'b0000000001000010   ;
13'd2167:weight<=16'b0000000001010010   ;
13'd2168:weight<=16'b0000000000000001   ;
13'd2169:weight<=16'b0000000010011110   ;
13'd2170:weight<=16'b1111111111100000   ;
13'd2171:weight<=16'b0000001000101000   ;
13'd2172:weight<=16'b1111111101111010   ;
13'd2173:weight<=16'b0000000101011101   ;
13'd2174:weight<=16'b0000010101111000   ;
13'd2175:weight<=16'b0000010100000110   ;
13'd2176:weight<=16'b1111101011010011   ;
13'd2177:weight<=16'b1111101001101101   ;
13'd2178:weight<=16'b1111110111010000   ;
13'd2179:weight<=16'b0000000100001111   ;
13'd2180:weight<=16'b1111111111011011   ;
13'd2181:weight<=16'b1111111110110110   ;
13'd2182:weight<=16'b0000000001011011   ;
13'd2183:weight<=16'b0000000100010011   ;
13'd2184:weight<=16'b1111111101011011   ;
13'd2185:weight<=16'b1111111111011001   ;
13'd2186:weight<=16'b0000000000100001   ;
13'd2187:weight<=16'b0000000001110100   ;
13'd2188:weight<=16'b0000000000001111   ;
13'd2189:weight<=16'b1111111110001010   ;
13'd2190:weight<=16'b1111111111000100   ;
13'd2191:weight<=16'b1111111111100111   ;
13'd2192:weight<=16'b1111111111100011   ;
13'd2193:weight<=16'b1111111110100101   ;
13'd2194:weight<=16'b0000000000100010   ;
13'd2195:weight<=16'b1111111111101111   ;
13'd2196:weight<=16'b0000000001000011   ;
13'd2197:weight<=16'b0000000001010000   ;
13'd2198:weight<=16'b1111111111100111   ;
13'd2199:weight<=16'b0000000001100011   ;
13'd2200:weight<=16'b0000000000110001   ;
13'd2201:weight<=16'b0000000000000101   ;
13'd2202:weight<=16'b0000000000010000   ;
13'd2203:weight<=16'b1111111110000000   ;
13'd2204:weight<=16'b1111111111100101   ;
13'd2205:weight<=16'b0000000011000010   ;
13'd2206:weight<=16'b1111111110011000   ;
13'd2207:weight<=16'b0000000001011010   ;
13'd2208:weight<=16'b0000000010001010   ;
13'd2209:weight<=16'b1111111100101011   ;
13'd2210:weight<=16'b1111111101100100   ;
13'd2211:weight<=16'b1111111110001111   ;
13'd2212:weight<=16'b1111111111000011   ;
13'd2213:weight<=16'b0000000000110110   ;
13'd2214:weight<=16'b1111111111100010   ;
13'd2215:weight<=16'b0000000000111011   ;
13'd2216:weight<=16'b0000000001000010   ;
13'd2217:weight<=16'b0000000001010010   ;
13'd2218:weight<=16'b0000000000000001   ;
13'd2219:weight<=16'b0000000010011110   ;
13'd2220:weight<=16'b1111111101101100   ;
13'd2221:weight<=16'b0000000000110000   ;
13'd2222:weight<=16'b0000000000011001   ;
13'd2223:weight<=16'b1111111101111011   ;
13'd2224:weight<=16'b1111111111001010   ;
13'd2225:weight<=16'b0000000000101011   ;
13'd2226:weight<=16'b0000000000010010   ;
13'd2227:weight<=16'b0000000000100101   ;
13'd2228:weight<=16'b0000000010100011   ;
13'd2229:weight<=16'b0000000000101000   ;
13'd2230:weight<=16'b1111111111011011   ;
13'd2231:weight<=16'b1111111110110110   ;
13'd2232:weight<=16'b0000000001011011   ;
13'd2233:weight<=16'b0000000100010011   ;
13'd2234:weight<=16'b1111111101011011   ;
13'd2235:weight<=16'b1111111111011001   ;
13'd2236:weight<=16'b0000000000100001   ;
13'd2237:weight<=16'b0000000001110100   ;
13'd2238:weight<=16'b0000000000001111   ;
13'd2239:weight<=16'b1111111110001010   ;
13'd2240:weight<=16'b1111111101001111   ;
13'd2241:weight<=16'b1111111100011010   ;
13'd2242:weight<=16'b0000000000011101   ;
13'd2243:weight<=16'b0000000100110110   ;
13'd2244:weight<=16'b0000000001011100   ;
13'd2245:weight<=16'b0000000000100000   ;
13'd2246:weight<=16'b1111111111011110   ;
13'd2247:weight<=16'b1111111100110010   ;
13'd2248:weight<=16'b0000000100100010   ;
13'd2249:weight<=16'b1111111110010101   ;
13'd2250:weight<=16'b0000000000110001   ;
13'd2251:weight<=16'b0000000000000101   ;
13'd2252:weight<=16'b0000000000010000   ;
13'd2253:weight<=16'b1111111110000000   ;
13'd2254:weight<=16'b1111111111100101   ;
13'd2255:weight<=16'b0000000011000010   ;
13'd2256:weight<=16'b1111111110011000  ;
13'd2257:weight<=16'b0000000001011010   ;
13'd2258:weight<=16'b0000000010001010   ;
13'd2259:weight<=16'b1111111100101011   ;
13'd2260:weight<=16'b0000000001001011   ;
13'd2261:weight<=16'b1111111111000111   ;
13'd2262:weight<=16'b0000000000011111   ;
13'd2263:weight<=16'b0000000000011001   ;
13'd2264:weight<=16'b0000000001010111   ;
13'd2265:weight<=16'b1111111111110111   ;
13'd2266:weight<=16'b1111111110101111   ;
13'd2267:weight<=16'b1111111111101100   ;
13'd2268:weight<=16'b1111111111011011   ;
13'd2269:weight<=16'b1111111111011010   ;
13'd2270:weight<=16'b1111111101101100   ;
13'd2271:weight<=16'b0000000000110000   ;
13'd2272:weight<=16'b0000000000011001   ;
13'd2273:weight<=16'b1111111101111011   ;
13'd2274:weight<=16'b1111111111001010   ;
13'd2275:weight<=16'b0000000000101011   ;
13'd2276:weight<=16'b0000000000010010   ;
13'd2277:weight<=16'b0000000000100101   ;
13'd2278:weight<=16'b0000000010100011   ;
13'd2279:weight<=16'b0000000000101000   ;
13'd2280:weight<=16'b1111111111000100   ;
13'd2281:weight<=16'b0000000110000011   ;
13'd2282:weight<=16'b1111111111110010   ;
13'd2283:weight<=16'b1111111100000101   ;
13'd2284:weight<=16'b1111111011011110   ;
13'd2285:weight<=16'b0000000011111101   ;
13'd2286:weight<=16'b1111111111101100   ;
13'd2287:weight<=16'b1111111111111010   ;
13'd2288:weight<=16'b0000000001011011   ;
13'd2289:weight<=16'b0000000000000101   ;
13'd2290:weight<=16'b1111111101001111   ;
13'd2291:weight<=16'b1111111100011010   ;
13'd2292:weight<=16'b0000000000011101   ;
13'd2293:weight<=16'b0000000100110110   ;
13'd2294:weight<=16'b0000000001011100   ;
13'd2295:weight<=16'b0000000000100000   ;
13'd2296:weight<=16'b1111111111011110   ;
13'd2297:weight<=16'b1111111100110010   ;
13'd2298:weight<=16'b0000000100100010   ;
13'd2299:weight<=16'b1111111110010101   ;
13'd2300:weight<=16'b0000000000001001   ;
13'd2301:weight<=16'b0000000000001100   ;
13'd2302:weight<=16'b0000000000000011   ;
13'd2303:weight<=16'b1111111110100000   ;
13'd2304:weight<=16'b0000000001111110   ;
13'd2305:weight<=16'b0000000000000000   ;
13'd2306:weight<=16'b1111111101111001   ;
13'd2307:weight<=16'b0000000001011001   ;
13'd2308:weight<=16'b1111111110100011   ;
13'd2309:weight<=16'b0000000010011000   ;
13'd2310:weight<=16'b0000000001001011   ;
13'd2311:weight<=16'b1111111111000111   ;
13'd2312:weight<=16'b0000000000011111   ;
13'd2313:weight<=16'b0000000000011001   ;
13'd2314:weight<=16'b0000000001010111   ;
13'd2315:weight<=16'b1111111111110111   ;
13'd2316:weight<=16'b1111111110101111   ;
13'd2317:weight<=16'b1111111111101100   ;
13'd2318:weight<=16'b1111111111011011   ;
13'd2319:weight<=16'b1111111111011010   ;
13'd2320:weight<=16'b1111111100111010   ;
13'd2321:weight<=16'b1111111111010100   ;
13'd2322:weight<=16'b1111111111010000   ;
13'd2323:weight<=16'b1111111101111010   ;
13'd2324:weight<=16'b1111111111100001   ;
13'd2325:weight<=16'b0000000111111001   ;
13'd2326:weight<=16'b0000000000111101   ;
13'd2327:weight<=16'b1111111111110001   ;
13'd2328:weight<=16'b1111111111101101   ;
13'd2329:weight<=16'b1111111111101000   ;
13'd2330:weight<=16'b1111111111000100   ;
13'd2331:weight<=16'b0000000110000011   ;
13'd2332:weight<=16'b1111111111110010   ;
13'd2333:weight<=16'b1111111100000101   ;
13'd2334:weight<=16'b1111111011011110   ;
13'd2335:weight<=16'b0000000011111101   ;
13'd2336:weight<=16'b1111111111101100   ;
13'd2337:weight<=16'b1111111111111010   ;
13'd2338:weight<=16'b0000000001011011   ;
13'd2339:weight<=16'b0000000000000101   ;
13'd2340:weight<=16'b1111111110101101   ;
13'd2341:weight<=16'b1111111110100100   ;
13'd2342:weight<=16'b1111111111111000   ;
13'd2343:weight<=16'b1111111111100001   ;
13'd2344:weight<=16'b1111111111001000   ;
13'd2345:weight<=16'b1111111111101111   ;
13'd2346:weight<=16'b0000000010100000   ;
13'd2347:weight<=16'b0000000000100001   ;
13'd2348:weight<=16'b0000000000111010   ;
13'd2349:weight<=16'b0000000000010111   ;
13'd2350:weight<=16'b0000000000001001   ;
13'd2351:weight<=16'b0000000000001100   ;
13'd2352:weight<=16'b0000000000000011   ;
13'd2353:weight<=16'b1111111110100000   ;
13'd2354:weight<=16'b0000000001111110   ;
13'd2355:weight<=16'b0000000000000000   ;
13'd2356:weight<=16'b1111111101111001   ;
13'd2357:weight<=16'b0000000001011001   ;
13'd2358:weight<=16'b1111111110100011   ;
13'd2359:weight<=16'b0000000010011000   ;
13'd2360:weight<=16'b1111111110111100   ;
13'd2361:weight<=16'b0000000001010000   ;
13'd2362:weight<=16'b0000000000001010   ;
13'd2363:weight<=16'b1111111101010001   ;
13'd2364:weight<=16'b0000000001011100   ;
13'd2365:weight<=16'b0000000010100110   ;
13'd2366:weight<=16'b1111111111011011   ;
13'd2367:weight<=16'b1111111100110110   ;
13'd2368:weight<=16'b0000000000111101   ;
13'd2369:weight<=16'b0000000010000000   ;
13'd2370:weight<=16'b1111111100111010   ;
13'd2371:weight<=16'b1111111111010100   ;
13'd2372:weight<=16'b1111111111010000   ;
13'd2373:weight<=16'b1111111101111010   ;
13'd2374:weight<=16'b1111111111100001   ;
13'd2375:weight<=16'b0000000111111001   ;
13'd2376:weight<=16'b0000000000111101   ;
13'd2377:weight<=16'b1111111111110001   ;
13'd2378:weight<=16'b1111111111101101   ;
13'd2379:weight<=16'b1111111111101000   ;
13'd2380:weight<=16'b0000000001100111   ;
13'd2381:weight<=16'b1111111110110000   ;
13'd2382:weight<=16'b1111111111000101   ;
13'd2383:weight<=16'b1111111111111111   ;
13'd2384:weight<=16'b1111111111111011   ;
13'd2385:weight<=16'b0000000001011111   ;
13'd2386:weight<=16'b0000000000111001   ;
13'd2387:weight<=16'b0000000000010101   ;
13'd2388:weight<=16'b0000000000111011   ;
13'd2389:weight<=16'b1111111101010001   ;
13'd2390:weight<=16'b1111111110101101   ;
13'd2391:weight<=16'b1111111110100100   ;
13'd2392:weight<=16'b1111111111111000   ;
13'd2393:weight<=16'b1111111111100001   ;
13'd2394:weight<=16'b1111111111001000   ;
13'd2395:weight<=16'b1111111111101111   ;
13'd2396:weight<=16'b0000000010100000   ;
13'd2397:weight<=16'b0000000000100001   ;
13'd2398:weight<=16'b0000000000111010   ;
13'd2399:weight<=16'b0000000000010111   ;
13'd2400:weight<=16'b0000000000101111   ;
13'd2401:weight<=16'b1111111111011000   ;
13'd2402:weight<=16'b1111111111001001   ;
13'd2403:weight<=16'b0000000000110001   ;
13'd2404:weight<=16'b1111111110110000   ;
13'd2405:weight<=16'b0000000001101101   ;
13'd2406:weight<=16'b1111111111110011   ;
13'd2407:weight<=16'b1111111110111010   ;
13'd2408:weight<=16'b0000000010010001   ;
13'd2409:weight<=16'b1111111110111001   ;
13'd2410:weight<=16'b1111111110111100   ;
13'd2411:weight<=16'b0000000001010000   ;
13'd2412:weight<=16'b0000000000001010   ;
13'd2413:weight<=16'b1111111101010001   ;
13'd2414:weight<=16'b0000000001011100   ;
13'd2415:weight<=16'b0000000010100110   ;
13'd2416:weight<=16'b1111111111011011   ;
13'd2417:weight<=16'b1111111100110110   ;
13'd2418:weight<=16'b0000000000111101   ;
13'd2419:weight<=16'b0000000010000000   ;
13'd2420:weight<=16'b1111111110010010   ;
13'd2421:weight<=16'b0000000000000111   ;
13'd2422:weight<=16'b0000000011110011   ;
13'd2423:weight<=16'b1111111111000000   ;
13'd2424:weight<=16'b1111111111010110   ;
13'd2425:weight<=16'b0000000000101000   ;
13'd2426:weight<=16'b0000000001000110   ;
13'd2427:weight<=16'b1111111111001011   ;
13'd2428:weight<=16'b1111111111100011   ;
13'd2429:weight<=16'b1111111111001101   ;
13'd2430:weight<=16'b0000000001100111   ;
13'd2431:weight<=16'b1111111110110000   ;
13'd2432:weight<=16'b1111111111000101   ;
13'd2433:weight<=16'b1111111111111111   ;
13'd2434:weight<=16'b1111111111111011   ;
13'd2435:weight<=16'b0000000001011111   ;
13'd2436:weight<=16'b0000000000111001   ;
13'd2437:weight<=16'b0000000000010101   ;
13'd2438:weight<=16'b0000000000111011   ;
13'd2439:weight<=16'b1111111101010001   ;
13'd2440:weight<=16'b0000000001100010   ;
13'd2441:weight<=16'b1111111111011111   ;
13'd2442:weight<=16'b0000000000001001  ;
13'd2443:weight<=16'b0000000001111100   ;
13'd2444:weight<=16'b1111111101101001   ;
13'd2445:weight<=16'b0000000010101010   ;
13'd2446:weight<=16'b1111111101110010   ;
13'd2447:weight<=16'b0000000001111011   ;
13'd2448:weight<=16'b1111111111011101   ;
13'd2449:weight<=16'b1111111110100100   ;
13'd2450:weight<=16'b0000000000101111   ;
13'd2451:weight<=16'b1111111111011000   ;
13'd2452:weight<=16'b1111111111001001   ;
13'd2453:weight<=16'b0000000000110001   ;
13'd2454:weight<=16'b1111111110110000   ;
13'd2455:weight<=16'b0000000001101101   ;
13'd2456:weight<=16'b1111111111110011   ;
13'd2457:weight<=16'b1111111110111010   ;
13'd2458:weight<=16'b0000000010010001   ;
13'd2459:weight<=16'b1111111110111001   ;
13'd2460:weight<=16'b0000000000010010   ;
13'd2461:weight<=16'b1111111110111100   ;
13'd2462:weight<=16'b1111111110101101   ;
13'd2463:weight<=16'b0000000000101000   ;
13'd2464:weight<=16'b1111111110010011   ;
13'd2465:weight<=16'b0000000001111110   ;
13'd2466:weight<=16'b1111111111100111   ;
13'd2467:weight<=16'b0000000010101101   ;
13'd2468:weight<=16'b1111111111101110   ;
13'd2469:weight<=16'b0000000001000111   ;
13'd2470:weight<=16'b1111111110010010   ;
13'd2471:weight<=16'b0000000000000111   ;
13'd2472:weight<=16'b0000000011110011   ;
13'd2473:weight<=16'b1111111111000000   ;
13'd2474:weight<=16'b1111111111010110   ;
13'd2475:weight<=16'b0000000000101000   ;
13'd2476:weight<=16'b0000000001000110   ;
13'd2477:weight<=16'b1111111111001011   ;
13'd2478:weight<=16'b1111111111100011   ;
13'd2479:weight<=16'b1111111111001101   ;
13'd2480:weight<=16'b0000000000111111   ;
13'd2481:weight<=16'b0000000001111001   ;
13'd2482:weight<=16'b0000000001000000   ;
13'd2483:weight<=16'b0000000000010110   ;
13'd2484:weight<=16'b1111111100111101   ;
13'd2485:weight<=16'b0000000001110111   ;
13'd2486:weight<=16'b1111111111111101   ;
13'd2487:weight<=16'b0000000000011101   ;
13'd2488:weight<=16'b1111111110100011   ;
13'd2489:weight<=16'b1111111110000100   ;
13'd2490:weight<=16'b0000000001100010   ;
13'd2491:weight<=16'b1111111111011111   ;
13'd2492:weight<=16'b0000000000001001   ;
13'd2493:weight<=16'b0000000001111100   ;
13'd2494:weight<=16'b1111111101101001   ;
13'd2495:weight<=16'b0000000010101010   ;
13'd2496:weight<=16'b1111111101110010   ;
13'd2497:weight<=16'b0000000001111011   ;
13'd2498:weight<=16'b1111111111011101   ;
13'd2499:weight<=16'b1111111110100100   ;
13'd2500:weight<=16'b1111111111101001   ;
13'd2501:weight<=16'b1111111111001110   ;
13'd2502:weight<=16'b0000000001111011   ;
13'd2503:weight<=16'b0000000000110110   ;
13'd2504:weight<=16'b1111111111111110   ;
13'd2505:weight<=16'b1111111111101011   ;
13'd2506:weight<=16'b0000000000001010   ;
13'd2507:weight<=16'b1111111111100011   ;
13'd2508:weight<=16'b1111111101111111   ;
13'd2509:weight<=16'b0000000001100100   ;
13'd2510:weight<=16'b0000000000010010   ;
13'd2511:weight<=16'b1111111110111100   ;
13'd2512:weight<=16'b1111111110101101   ;
13'd2513:weight<=16'b0000000000101000   ;
13'd2514:weight<=16'b1111111110010011   ;
13'd2515:weight<=16'b0000000001111110   ;
13'd2516:weight<=16'b1111111111100111   ;
13'd2517:weight<=16'b0000000010101101   ;
13'd2518:weight<=16'b1111111111101110   ;
13'd2519:weight<=16'b0000000001000111   ;
13'd2520:weight<=16'b1111111111011110   ;
13'd2521:weight<=16'b0000000000100111   ;
13'd2522:weight<=16'b1111111111110100   ;
13'd2523:weight<=16'b0000000010111110   ;
13'd2524:weight<=16'b0000000000110111   ;
13'd2525:weight<=16'b1111111110110011   ;
13'd2526:weight<=16'b1111111111111011   ;
13'd2527:weight<=16'b0000000000100110   ;
13'd2528:weight<=16'b0000000000001000   ;
13'd2529:weight<=16'b1111111101110001   ;
13'd2530:weight<=16'b0000000000111111   ;
13'd2531:weight<=16'b0000000001111001   ;
13'd2532:weight<=16'b0000000001000000   ;
13'd2533:weight<=16'b0000000000010110   ;
13'd2534:weight<=16'b1111111100111101   ;
13'd2535:weight<=16'b0000000001110111   ;
13'd2536:weight<=16'b1111111111111101   ;
13'd2537:weight<=16'b0000000000011101   ;
13'd2538:weight<=16'b1111111110100011   ;
13'd2539:weight<=16'b1111111110000100   ;
13'd2540:weight<=16'b1111111110000011   ;
13'd2541:weight<=16'b1111111111000100   ;
13'd2542:weight<=16'b0000000010101101   ;
13'd2543:weight<=16'b1111111110011001   ;
13'd2544:weight<=16'b0000000010100011   ;
13'd2545:weight<=16'b1111111111100001   ;
13'd2546:weight<=16'b1111111110110110   ;
13'd2547:weight<=16'b1111111111000111   ;
13'd2548:weight<=16'b0000000001101100   ;
13'd2549:weight<=16'b0000000000011000   ;
13'd2550:weight<=16'b1111111111101001   ;
13'd2551:weight<=16'b1111111111001110   ;
13'd2552:weight<=16'b0000000001111011   ;
13'd2553:weight<=16'b0000000000110110   ;
13'd2554:weight<=16'b1111111111111110   ;
13'd2555:weight<=16'b1111111111101011   ;
13'd2556:weight<=16'b0000000000001010   ;
13'd2557:weight<=16'b1111111111100011   ;
13'd2558:weight<=16'b1111111101111111   ;
13'd2559:weight<=16'b0000000001100100   ;
13'd2560:weight<=16'b1111111110111001   ;
13'd2561:weight<=16'b1111111110011101   ;
13'd2562:weight<=16'b0000000000101000   ;
13'd2563:weight<=16'b1111111111010101   ;
13'd2564:weight<=16'b0000000111000100   ;
13'd2565:weight<=16'b1111111111110111   ;
13'd2566:weight<=16'b1111111111001010   ;
13'd2567:weight<=16'b0000000000111011   ;
13'd2568:weight<=16'b1111111100010110   ;
13'd2569:weight<=16'b1111111111111011   ;
13'd2570:weight<=16'b1111111111011110   ;
13'd2571:weight<=16'b0000000000100111   ;
13'd2572:weight<=16'b1111111111110100   ;
13'd2573:weight<=16'b0000000010111110   ;
13'd2574:weight<=16'b0000000000110111   ;
13'd2575:weight<=16'b1111111110110011   ;
13'd2576:weight<=16'b1111111111111011   ;
13'd2577:weight<=16'b0000000000100110   ;
13'd2578:weight<=16'b0000000000001000   ;
13'd2579:weight<=16'b1111111101110001   ;
13'd2580:weight<=16'b0000000001110001   ;
13'd2581:weight<=16'b1111111110100001   ;
13'd2582:weight<=16'b0000000001001100   ;
13'd2583:weight<=16'b1111111111010010   ;
13'd2584:weight<=16'b0000000011100111   ;
13'd2585:weight<=16'b1111111110000111   ;
13'd2586:weight<=16'b1111111111100100   ;
13'd2587:weight<=16'b0000000010110010   ;
13'd2588:weight<=16'b1111111011100110   ;
13'd2589:weight<=16'b0000000000011100   ;
13'd2590:weight<=16'b1111111110000011   ;
13'd2591:weight<=16'b1111111111000100   ;
13'd2592:weight<=16'b0000000010101101   ;
13'd2593:weight<=16'b1111111110011001   ;
13'd2594:weight<=16'b0000000010100011   ;
13'd2595:weight<=16'b1111111111100001   ;
13'd2596:weight<=16'b1111111110110110   ;
13'd2597:weight<=16'b1111111111000111   ;
13'd2598:weight<=16'b0000000001101100   ;
13'd2599:weight<=16'b0000000000011000   ;
13'd2600:weight<=16'b0000000000111011   ;
13'd2601:weight<=16'b1111111110100101   ;
13'd2602:weight<=16'b1111111111111000   ;
13'd2603:weight<=16'b0000000001100100   ;
13'd2604:weight<=16'b0000000000111001   ;
13'd2605:weight<=16'b0000000010110100   ;
13'd2606:weight<=16'b1111111110000010   ;
13'd2607:weight<=16'b1111111110100100   ;
13'd2608:weight<=16'b1111111111101100   ;
13'd2609:weight<=16'b1111111111101110   ;
13'd2610:weight<=16'b1111111110111001   ;
13'd2611:weight<=16'b1111111110011101   ;
13'd2612:weight<=16'b0000000000101000   ;
13'd2613:weight<=16'b1111111111010101   ;
13'd2614:weight<=16'b0000000111000100   ;
13'd2615:weight<=16'b1111111111110111   ;
13'd2616:weight<=16'b1111111111001010   ;
13'd2617:weight<=16'b0000000000111011   ;
13'd2618:weight<=16'b1111111100010110   ;
13'd2619:weight<=16'b1111111111111011   ;
13'd2620:weight<=16'b0000000000000011   ;
13'd2621:weight<=16'b0000000000011000   ;
13'd2622:weight<=16'b1111111111111011   ;
13'd2623:weight<=16'b1111111111100011   ;
13'd2624:weight<=16'b0000000000001001   ;
13'd2625:weight<=16'b0000000000001001   ;
13'd2626:weight<=16'b0000000000110000   ;
13'd2627:weight<=16'b1111111110011110   ;
13'd2628:weight<=16'b0000000000001011   ;
13'd2629:weight<=16'b0000000000101100   ;
13'd2630:weight<=16'b0000000001110001   ;
13'd2631:weight<=16'b1111111110100001   ;
13'd2632:weight<=16'b0000000001001100   ;
13'd2633:weight<=16'b1111111111010010   ;
13'd2634:weight<=16'b0000000011100111   ;
13'd2635:weight<=16'b1111111110000111   ;
13'd2636:weight<=16'b1111111111100100   ;
13'd2637:weight<=16'b0000000010110010   ;
13'd2638:weight<=16'b1111111011100110   ;
13'd2639:weight<=16'b0000000000011100   ;
13'd2640:weight<=16'b1111111110101010   ;
13'd2641:weight<=16'b0000000001001110   ;
13'd2642:weight<=16'b0000000000011001   ;
13'd2643:weight<=16'b0000000000110110   ;
13'd2644:weight<=16'b1111111111001111   ;
13'd2645:weight<=16'b1111111011111001   ;
13'd2646:weight<=16'b0000000001100100   ;
13'd2647:weight<=16'b0000000001001101   ;
13'd2648:weight<=16'b1111111111101110   ;
13'd2649:weight<=16'b0000000001110001   ;
13'd2650:weight<=16'b0000000000111011   ;
13'd2651:weight<=16'b1111111110100101   ;
13'd2652:weight<=16'b1111111111111000   ;
13'd2653:weight<=16'b0000000001100100   ;
13'd2654:weight<=16'b0000000000111001   ;
13'd2655:weight<=16'b0000000010110100   ;
13'd2656:weight<=16'b1111111110000010   ;
13'd2657:weight<=16'b1111111110100100   ;
13'd2658:weight<=16'b1111111111101100   ;
13'd2659:weight<=16'b1111111111101110   ;
13'd2660:weight<=16'b0000000000111111   ;
13'd2661:weight<=16'b1111111100100111   ;
13'd2662:weight<=16'b0000000000110100   ;
13'd2663:weight<=16'b1111111101110101   ;
13'd2664:weight<=16'b0000000000010101   ;
13'd2665:weight<=16'b0000000000111001   ;
13'd2666:weight<=16'b1111111111110011   ;
13'd2667:weight<=16'b0000000000001010   ;
13'd2668:weight<=16'b0000000000101100   ;
13'd2669:weight<=16'b0000000010000011   ;
13'd2670:weight<=16'b0000000000000011   ;
13'd2671:weight<=16'b0000000000011000   ;
13'd2672:weight<=16'b1111111111111011   ;
13'd2673:weight<=16'b1111111111100011   ;
13'd2674:weight<=16'b0000000000001001   ;
13'd2675:weight<=16'b0000000000001001   ;
13'd2676:weight<=16'b0000000000110000   ;
13'd2677:weight<=16'b1111111110011110   ;
13'd2678:weight<=16'b0000000000001011   ;
13'd2679:weight<=16'b0000000000101100   ;
13'd2680:weight<=16'b1111111111000101   ;
13'd2681:weight<=16'b0000000010000010   ;
13'd2682:weight<=16'b0000000000000110   ;
13'd2683:weight<=16'b1111111111001111   ;
13'd2684:weight<=16'b1111111110011011   ;
13'd2685:weight<=16'b0000000000011110  ;
13'd2686:weight<=16'b1111111110111011   ;
13'd2687:weight<=16'b0000000000010001   ;
13'd2688:weight<=16'b0000000100100100   ;
13'd2689:weight<=16'b1111111101010101   ;
13'd2690:weight<=16'b1111111110101010   ;
13'd2691:weight<=16'b0000000001001110   ;
13'd2692:weight<=16'b0000000000011001   ;
13'd2693:weight<=16'b0000000000110110   ;
13'd2694:weight<=16'b1111111111001111   ;
13'd2695:weight<=16'b1111111011111001   ;
13'd2696:weight<=16'b0000000001100100   ;
13'd2697:weight<=16'b0000000001001101   ;
13'd2698:weight<=16'b1111111111101110   ;
13'd2699:weight<=16'b0000000001110001   ;
13'd2700:weight<=16'b0000000000011001   ;
13'd2701:weight<=16'b1111111111010101   ;
13'd2702:weight<=16'b1111111111011011   ;
13'd2703:weight<=16'b0000000010011111   ;
13'd2704:weight<=16'b1111111101011011   ;
13'd2705:weight<=16'b1111111111110110   ;
13'd2706:weight<=16'b0000000001100010   ;
13'd2707:weight<=16'b1111111111001010   ;
13'd2708:weight<=16'b0000000001111101   ;
13'd2709:weight<=16'b1111111111001111   ;
13'd2710:weight<=16'b0000000000111111   ;
13'd2711:weight<=16'b1111111100100111   ;
13'd2712:weight<=16'b0000000000110100   ;
13'd2713:weight<=16'b1111111101110101   ;
13'd2714:weight<=16'b0000000000010101   ;
13'd2715:weight<=16'b0000000000111001   ;
13'd2716:weight<=16'b1111111111110011   ;
13'd2717:weight<=16'b0000000000001010   ;
13'd2718:weight<=16'b0000000000101100   ;
13'd2719:weight<=16'b0000000010000011   ;
13'd2720:weight<=16'b1111111101101100   ;
13'd2721:weight<=16'b0000000001011000   ;
13'd2722:weight<=16'b0000000101010000   ;
13'd2723:weight<=16'b0000000011000000   ;
13'd2724:weight<=16'b0000000110111111   ;
13'd2725:weight<=16'b0000000001000110   ;
13'd2726:weight<=16'b1111111100010100   ;
13'd2727:weight<=16'b1111111010001101   ;
13'd2728:weight<=16'b1111111111110010   ;
13'd2729:weight<=16'b1111111100010000   ;
13'd2730:weight<=16'b1111111111000101   ;
13'd2731:weight<=16'b0000000010000010   ;
13'd2732:weight<=16'b0000000000000110   ;
13'd2733:weight<=16'b1111111111001111   ;
13'd2734:weight<=16'b1111111110011011   ;
13'd2735:weight<=16'b0000000000011110   ;
13'd2736:weight<=16'b1111111110111011   ;
13'd2737:weight<=16'b0000000000010001   ;
13'd2738:weight<=16'b0000000100100100   ;
13'd2739:weight<=16'b1111111101010101   ;
13'd2740:weight<=16'b1111111111111110   ;
13'd2741:weight<=16'b1111111110001100   ;
13'd2742:weight<=16'b0000000011010000   ;
13'd2743:weight<=16'b0000000000001110   ;
13'd2744:weight<=16'b0000000000000100   ;
13'd2745:weight<=16'b1111111111001001   ;
13'd2746:weight<=16'b1111111111101011   ;
13'd2747:weight<=16'b1111111111111100   ;
13'd2748:weight<=16'b1111111111101101   ;
13'd2749:weight<=16'b1111111111101101   ;
13'd2750:weight<=16'b0000000000011001   ;
13'd2751:weight<=16'b1111111111010101   ;
13'd2752:weight<=16'b1111111111011011   ;
13'd2753:weight<=16'b0000000010011111   ;
13'd2754:weight<=16'b1111111101011011   ;
13'd2755:weight<=16'b1111111111110110   ;
13'd2756:weight<=16'b0000000001100010   ;
13'd2757:weight<=16'b1111111111001010   ;
13'd2758:weight<=16'b0000000001111101   ;
13'd2759:weight<=16'b1111111111001111   ;
13'd2760:weight<=16'b0000000001010101   ;
13'd2761:weight<=16'b0000000001011010   ;
13'd2762:weight<=16'b1111111111100001   ;
13'd2763:weight<=16'b0000000001111011   ;
13'd2764:weight<=16'b1111111110110000   ;
13'd2765:weight<=16'b1111111101100011   ;
13'd2766:weight<=16'b1111111111110011   ;
13'd2767:weight<=16'b1111111111010000   ;
13'd2768:weight<=16'b0000000000100010   ;
13'd2769:weight<=16'b0000000001010110   ;
13'd2770:weight<=16'b1111111101101100   ;
13'd2771:weight<=16'b0000000001011000   ;
13'd2772:weight<=16'b0000000101010000   ;
13'd2773:weight<=16'b0000000011000000   ;
13'd2774:weight<=16'b0000000110111111   ;
13'd2775:weight<=16'b0000000001000110   ;
13'd2776:weight<=16'b1111111100010100   ;
13'd2777:weight<=16'b1111111010001101   ;
13'd2778:weight<=16'b1111111111110010   ;
13'd2779:weight<=16'b1111111100010000   ;
13'd2780:weight<=16'b1111111111100101   ;
13'd2781:weight<=16'b1111111100101100   ;
13'd2782:weight<=16'b0000001000000100   ;
13'd2783:weight<=16'b0000000001110110   ;
13'd2784:weight<=16'b0000000010000001   ;
13'd2785:weight<=16'b1111111111101100   ;
13'd2786:weight<=16'b1111111101101001   ;
13'd2787:weight<=16'b1111111011000111   ;
13'd2788:weight<=16'b1111111111011001   ;
13'd2789:weight<=16'b0000000000011100   ;
13'd2790:weight<=16'b1111111111111110   ;
13'd2791:weight<=16'b1111111110001100   ;
13'd2792:weight<=16'b0000000011010000   ;
13'd2793:weight<=16'b0000000000001110   ;
13'd2794:weight<=16'b0000000000000100   ;
13'd2795:weight<=16'b1111111111001001   ;
13'd2796:weight<=16'b1111111111101011   ;
13'd2797:weight<=16'b1111111111111100   ;
13'd2798:weight<=16'b1111111111101101   ;
13'd2799:weight<=16'b1111111111101101   ;
13'd2800:weight<=16'b0000000001100000   ;
13'd2801:weight<=16'b1111111111000111   ;
13'd2802:weight<=16'b1111111100000100   ;
13'd2803:weight<=16'b1111111111010001   ;
13'd2804:weight<=16'b1111111111010000   ;
13'd2805:weight<=16'b0000000000101011   ;
13'd2806:weight<=16'b0000000001010000   ;
13'd2807:weight<=16'b0000000001011110   ;
13'd2808:weight<=16'b0000000000110110   ;
13'd2809:weight<=16'b0000000001001011   ;
13'd2810:weight<=16'b0000000001010101   ;
13'd2811:weight<=16'b0000000001011010   ;
13'd2812:weight<=16'b1111111111100001   ;
13'd2813:weight<=16'b0000000001111011   ;
13'd2814:weight<=16'b1111111110110000   ;
13'd2815:weight<=16'b1111111101100011   ;
13'd2816:weight<=16'b1111111111110011   ;
13'd2817:weight<=16'b1111111111010000   ;
13'd2818:weight<=16'b0000000000100010   ;
13'd2819:weight<=16'b0000000001010110   ;
13'd2820:weight<=16'b1111111111011100   ;
13'd2821:weight<=16'b1111111111100000   ;
13'd2822:weight<=16'b1111111101100111   ;
13'd2823:weight<=16'b0000000000000100   ;
13'd2824:weight<=16'b0000000000101100   ;
13'd2825:weight<=16'b0000000000110000   ;
13'd2826:weight<=16'b0000000001100011   ;
13'd2827:weight<=16'b0000000000110011   ;
13'd2828:weight<=16'b1111111111011110   ;
13'd2829:weight<=16'b0000000000011111   ;
13'd2830:weight<=16'b1111111111100101   ;
13'd2831:weight<=16'b1111111100101100   ;
13'd2832:weight<=16'b0000001000000100   ;
13'd2833:weight<=16'b0000000001110110   ;
13'd2834:weight<=16'b0000000010000001   ;
13'd2835:weight<=16'b1111111111101100   ;
13'd2836:weight<=16'b1111111101101001   ;
13'd2837:weight<=16'b1111111011000111   ;
13'd2838:weight<=16'b1111111111011001   ;
13'd2839:weight<=16'b0000000000011100   ;
13'd2840:weight<=16'b0000000001001111   ;
13'd2841:weight<=16'b1111111110111101   ;
13'd2842:weight<=16'b1111111111100000   ;
13'd2843:weight<=16'b1111111111010111   ;
13'd2844:weight<=16'b0000000000100101   ;
13'd2845:weight<=16'b0000000000011101   ;
13'd2846:weight<=16'b0000000000100011   ;
13'd2847:weight<=16'b0000000001101001   ;
13'd2848:weight<=16'b1111111101111100   ;
13'd2849:weight<=16'b1111111111111011   ;
13'd2850:weight<=16'b0000000001100000   ;
13'd2851:weight<=16'b1111111111000111   ;
13'd2852:weight<=16'b1111111100000100   ;
13'd2853:weight<=16'b1111111111010001   ;
13'd2854:weight<=16'b1111111111010000   ;
13'd2855:weight<=16'b0000000000101011   ;
13'd2856:weight<=16'b0000000001010000   ;
13'd2857:weight<=16'b0000000001011110   ;
13'd2858:weight<=16'b0000000000110110   ;
13'd2859:weight<=16'b0000000001001011   ;
13'd2860:weight<=16'b1111111101011111   ;
13'd2861:weight<=16'b0000000000000000   ;
13'd2862:weight<=16'b0000000000000010   ;
13'd2863:weight<=16'b1111111111010001   ;
13'd2864:weight<=16'b0000000101000101   ;
13'd2865:weight<=16'b1111111111010111   ;
13'd2866:weight<=16'b1111111110001010   ;
13'd2867:weight<=16'b1111111110110011   ;
13'd2868:weight<=16'b0000000011000100   ;
13'd2869:weight<=16'b1111111111000101   ;
13'd2870:weight<=16'b1111111111011100   ;
13'd2871:weight<=16'b1111111111100000   ;
13'd2872:weight<=16'b1111111101100111   ;
13'd2873:weight<=16'b0000000000000100   ;
13'd2874:weight<=16'b0000000000101100   ;
13'd2875:weight<=16'b0000000000110000   ;
13'd2876:weight<=16'b0000000001100011   ;
13'd2877:weight<=16'b0000000000110011   ;
13'd2878:weight<=16'b1111111111011110   ;
13'd2879:weight<=16'b0000000000011111   ;
13'd2880:weight<=16'b0000000010011110   ;
13'd2881:weight<=16'b1111111101110000   ;
13'd2882:weight<=16'b0000000100111110   ;
13'd2883:weight<=16'b0000000101110110   ;
13'd2884:weight<=16'b1111111101001001   ;
13'd2885:weight<=16'b1111110110110101   ;
13'd2886:weight<=16'b1111110111010110   ;
13'd2887:weight<=16'b0000000011100001   ;
13'd2888:weight<=16'b0000000000100100   ;
13'd2889:weight<=16'b0000000110011001   ;
13'd2890:weight<=16'b0000000001001111   ;
13'd2891:weight<=16'b1111111110111101   ;
13'd2892:weight<=16'b1111111111100000   ;
13'd2893:weight<=16'b1111111111010111   ;
13'd2894:weight<=16'b0000000000100101   ;
13'd2895:weight<=16'b0000000000011101   ;
13'd2896:weight<=16'b0000000000100011   ;
13'd2897:weight<=16'b0000000001101001   ;
13'd2898:weight<=16'b1111111101111100   ;
13'd2899:weight<=16'b1111111111111011   ;
13'd2900:weight<=16'b0000000000010110   ;
13'd2901:weight<=16'b0000000001001000   ;
13'd2902:weight<=16'b1111111110001111   ;
13'd2903:weight<=16'b1111111101101101   ;
13'd2904:weight<=16'b1111111110011000   ;
13'd2905:weight<=16'b0000000010010100   ;
13'd2906:weight<=16'b1111111111000100   ;
13'd2907:weight<=16'b1111111111011101   ;
13'd2908:weight<=16'b0000000001001111   ;
13'd2909:weight<=16'b0000000011001000   ;
13'd2910:weight<=16'b1111111101011111   ;
13'd2911:weight<=16'b0000000000000000   ;
13'd2912:weight<=16'b0000000000000010   ;
13'd2913:weight<=16'b1111111111010001   ;
13'd2914:weight<=16'b0000000101000101   ;
13'd2915:weight<=16'b1111111111010111   ;
13'd2916:weight<=16'b1111111110001010   ;
13'd2917:weight<=16'b1111111110110011   ;
13'd2918:weight<=16'b0000000011000100   ;
13'd2919:weight<=16'b1111111111000101   ;
13'd2920:weight<=16'b1111111101100101   ;
13'd2921:weight<=16'b1111111101100111   ;
13'd2922:weight<=16'b0000000001110101   ;
13'd2923:weight<=16'b1111111011111101   ;
13'd2924:weight<=16'b0000000001010110   ;
13'd2925:weight<=16'b0000000000010111   ;
13'd2926:weight<=16'b1111111110010111   ;
13'd2927:weight<=16'b0000000010011110   ;
13'd2928:weight<=16'b0000000010101001   ;
13'd2929:weight<=16'b0000000010111100   ;
13'd2930:weight<=16'b0000000010011110   ;
13'd2931:weight<=16'b1111111101110000   ;
13'd2932:weight<=16'b0000000100111110   ;
13'd2933:weight<=16'b0000000101110110   ;
13'd2934:weight<=16'b1111111101001001   ;
13'd2935:weight<=16'b1111110110110101   ;
13'd2936:weight<=16'b1111110111010110   ;
13'd2937:weight<=16'b0000000011100001   ;
13'd2938:weight<=16'b0000000000100100   ;
13'd2939:weight<=16'b0000000110011001   ;
13'd2940:weight<=16'b1111111111100000   ;
13'd2941:weight<=16'b1111111111000000   ;
13'd2942:weight<=16'b0000000101110000   ;
13'd2943:weight<=16'b0000000000010100   ;
13'd2944:weight<=16'b0000000010010100   ;
13'd2945:weight<=16'b1111111110011101   ;
13'd2946:weight<=16'b1111111100101110   ;
13'd2947:weight<=16'b1111111111011010   ;
13'd2948:weight<=16'b1111111111010000   ;
13'd2949:weight<=16'b1111111111111001   ;
13'd2950:weight<=16'b0000000000010110   ;
13'd2951:weight<=16'b0000000001001000   ;
13'd2952:weight<=16'b1111111110001111   ;
13'd2953:weight<=16'b1111111101101101   ;
13'd2954:weight<=16'b1111111110011000   ;
13'd2955:weight<=16'b0000000010010100   ;
13'd2956:weight<=16'b1111111111000100   ;
13'd2957:weight<=16'b1111111111011101   ;
13'd2958:weight<=16'b0000000001001111   ;
13'd2959:weight<=16'b0000000011001000   ;
13'd2960:weight<=16'b0000000100011010   ;
13'd2961:weight<=16'b0000000001110010   ;
13'd2962:weight<=16'b1111111110000010   ;
13'd2963:weight<=16'b1111111111110110   ;
13'd2964:weight<=16'b0000000001110010   ;
13'd2965:weight<=16'b1111111110110101   ;
13'd2966:weight<=16'b1111111100010000   ;
13'd2967:weight<=16'b0000000100001001   ;
13'd2968:weight<=16'b0000000000010010   ;
13'd2969:weight<=16'b1111111100010100   ;
13'd2970:weight<=16'b1111111101100101   ;
13'd2971:weight<=16'b1111111101100111   ;
13'd2972:weight<=16'b0000000001110101   ;
13'd2973:weight<=16'b1111111011111101   ;
13'd2974:weight<=16'b0000000001010110   ;
13'd2975:weight<=16'b0000000000010111   ;
13'd2976:weight<=16'b1111111110010111   ;
13'd2977:weight<=16'b0000000010011110   ;
13'd2978:weight<=16'b0000000010101001   ;
13'd2979:weight<=16'b0000000010111100   ;
13'd2980:weight<=16'b1111111111001111   ;
13'd2981:weight<=16'b1111111110111001   ;
13'd2982:weight<=16'b0000000000011000   ;
13'd2983:weight<=16'b1111111110110011   ;
13'd2984:weight<=16'b0000000000001100   ;
13'd2985:weight<=16'b0000000010011100   ;
13'd2986:weight<=16'b1111111111000010   ;
13'd2987:weight<=16'b0000000000100011   ;
13'd2988:weight<=16'b0000000001101001   ;
13'd2989:weight<=16'b1111111111001010   ;
13'd2990:weight<=16'b1111111111100000   ;
13'd2991:weight<=16'b1111111111000000   ;
13'd2992:weight<=16'b0000000101110000   ;
13'd2993:weight<=16'b0000000000010100   ;
13'd2994:weight<=16'b0000000010010100   ;
13'd2995:weight<=16'b1111111110011101   ;
13'd2996:weight<=16'b1111111100101110   ;
13'd2997:weight<=16'b1111111111011010   ;
13'd2998:weight<=16'b1111111111010000   ;
13'd2999:weight<=16'b1111111111111001   ;
13'd3000:weight<=16'b0000000000100100   ;
13'd3001:weight<=16'b0000000001101010   ;
13'd3002:weight<=16'b1111111111111110   ;
13'd3003:weight<=16'b1111111111001110   ;
13'd3004:weight<=16'b0000000010011000   ;
13'd3005:weight<=16'b0000000000111010   ;
13'd3006:weight<=16'b1111111111000110   ;
13'd3007:weight<=16'b1111111111100000   ;
13'd3008:weight<=16'b1111111111000001   ;
13'd3009:weight<=16'b1111111110101110   ;
13'd3010:weight<=16'b0000000100011010   ;
13'd3011:weight<=16'b0000000001110010   ;
13'd3012:weight<=16'b1111111110000010   ;
13'd3013:weight<=16'b1111111111110110   ;
13'd3014:weight<=16'b0000000001110010   ;
13'd3015:weight<=16'b1111111110110101   ;
13'd3016:weight<=16'b1111111100010000   ;
13'd3017:weight<=16'b0000000100001001   ;
13'd3018:weight<=16'b0000000000010010   ;
13'd3019:weight<=16'b1111111100010100   ;
13'd3020:weight<=16'b1111111111110101   ;
13'd3021:weight<=16'b0000000001101010   ;
13'd3022:weight<=16'b0000000011110010   ;
13'd3023:weight<=16'b1111111111000000   ;
13'd3024:weight<=16'b1111111111110110   ;
13'd3025:weight<=16'b0000000010011001   ;
13'd3026:weight<=16'b1111111111111101   ;
13'd3027:weight<=16'b1111111110100010   ;
13'd3028:weight<=16'b1111111100010110   ;
13'd3029:weight<=16'b1111111111100101   ;
13'd3030:weight<=16'b1111111111001111   ;
13'd3031:weight<=16'b1111111110111001   ;
13'd3032:weight<=16'b0000000000011000   ;
13'd3033:weight<=16'b1111111110110011   ;
13'd3034:weight<=16'b0000000000001100   ;
13'd3035:weight<=16'b0000000010011100   ;
13'd3036:weight<=16'b1111111111000010   ;
13'd3037:weight<=16'b0000000000100011   ;
13'd3038:weight<=16'b0000000001101001   ;
13'd3039:weight<=16'b1111111111001010   ;
13'd3040:weight<=16'b1111111100100101   ;
13'd3041:weight<=16'b0000000000000111   ;
13'd3042:weight<=16'b0000000001101100   ;
13'd3043:weight<=16'b1111111101110100   ;
13'd3044:weight<=16'b0000000010010100   ;
13'd3045:weight<=16'b0000000100000101   ;
13'd3046:weight<=16'b1111111100110010   ;
13'd3047:weight<=16'b0000000100111101   ;
13'd3048:weight<=16'b1111111111111011   ;
13'd3049:weight<=16'b1111111110010010   ;
13'd3050:weight<=16'b0000000000100100   ;
13'd3051:weight<=16'b0000000001101010   ;
13'd3052:weight<=16'b1111111111111110   ;
13'd3053:weight<=16'b1111111111001110   ;
13'd3054:weight<=16'b0000000010011000   ;
13'd3055:weight<=16'b0000000000111010   ;
13'd3056:weight<=16'b1111111111000110   ;
13'd3057:weight<=16'b1111111111100000   ;
13'd3058:weight<=16'b1111111111000001   ;
13'd3059:weight<=16'b1111111110101110   ;
13'd3060:weight<=16'b1111111110010010   ;
13'd3061:weight<=16'b0000000001110010   ;
13'd3062:weight<=16'b1111111111111111   ;
13'd3063:weight<=16'b1111111111111001   ;
13'd3064:weight<=16'b0000000000000001   ;
13'd3065:weight<=16'b0000000000000000   ;
13'd3066:weight<=16'b1111111111010011   ;
13'd3067:weight<=16'b0000000000101010   ;
13'd3068:weight<=16'b0000000000000111   ;
13'd3069:weight<=16'b0000000000100000   ;
13'd3070:weight<=16'b1111111111110101   ;
13'd3071:weight<=16'b0000000001101010   ;
13'd3072:weight<=16'b0000000011110010   ;
13'd3073:weight<=16'b1111111111000000   ;
13'd3074:weight<=16'b1111111111110110   ;
13'd3075:weight<=16'b0000000010011001   ;
13'd3076:weight<=16'b1111111111111101   ;
13'd3077:weight<=16'b1111111110100010   ;
13'd3078:weight<=16'b1111111100010110   ;
13'd3079:weight<=16'b1111111111100101   ;
13'd3080:weight<=16'b1111111111101001   ;
13'd3081:weight<=16'b0000000001000111   ;
13'd3082:weight<=16'b1111111111001100   ;
13'd3083:weight<=16'b0000000000101101   ;
13'd3084:weight<=16'b0000000001110010   ;
13'd3085:weight<=16'b1111111110101101   ;
13'd3086:weight<=16'b0000000001111001   ;
13'd3087:weight<=16'b0000000001000110   ;
13'd3088:weight<=16'b1111111100100110   ;
13'd3089:weight<=16'b0000000000000011   ;
13'd3090:weight<=16'b1111111100100101  ;
13'd3091:weight<=16'b0000000000000111   ;
13'd3092:weight<=16'b0000000001101100   ;
13'd3093:weight<=16'b1111111101110100   ;
13'd3094:weight<=16'b0000000010010100   ;
13'd3095:weight<=16'b0000000100000101   ;
13'd3096:weight<=16'b1111111100110010   ;
13'd3097:weight<=16'b0000000100111101   ;
13'd3098:weight<=16'b1111111111111011   ;
13'd3099:weight<=16'b1111111110010010   ;
13'd3100:weight<=16'b1111111111111011   ;
13'd3101:weight<=16'b1111111101100000   ;
13'd3102:weight<=16'b0000000000111010   ;
13'd3103:weight<=16'b0000000001110011   ;
13'd3104:weight<=16'b0000000011110001   ;
13'd3105:weight<=16'b1111111110101000   ;
13'd3106:weight<=16'b0000000001100000   ;
13'd3107:weight<=16'b1111111110011111   ;
13'd3108:weight<=16'b1111111101001101   ;
13'd3109:weight<=16'b0000000001000000   ;
13'd3110:weight<=16'b1111111110010010   ;
13'd3111:weight<=16'b0000000001110010   ;
13'd3112:weight<=16'b1111111111111111   ;
13'd3113:weight<=16'b1111111111111001   ;
13'd3114:weight<=16'b0000000000000001   ;
13'd3115:weight<=16'b0000000000000000   ;
13'd3116:weight<=16'b1111111111010011   ;
13'd3117:weight<=16'b0000000000101010   ;
13'd3118:weight<=16'b0000000000000111   ;
13'd3119:weight<=16'b0000000000100000   ;
13'd3120:weight<=16'b1111111111101010   ;
13'd3121:weight<=16'b0000000001010010   ;
13'd3122:weight<=16'b0000000001010001   ;
13'd3123:weight<=16'b1111111101011100   ;
13'd3124:weight<=16'b0000000010110100   ;
13'd3125:weight<=16'b0000000010101011   ;
13'd3126:weight<=16'b1111111110110001   ;
13'd3127:weight<=16'b1111111101101000   ;
13'd3128:weight<=16'b1111111111000100   ;
13'd3129:weight<=16'b0000000000000001   ;
13'd3130:weight<=16'b1111111111101001   ;
13'd3131:weight<=16'b0000000001000111   ;
13'd3132:weight<=16'b1111111111001100   ;
13'd3133:weight<=16'b0000000000101101   ;
13'd3134:weight<=16'b0000000001110010   ;
13'd3135:weight<=16'b1111111110101101   ;
13'd3136:weight<=16'b0000000001111001   ;
13'd3137:weight<=16'b0000000001000110   ;
13'd3138:weight<=16'b1111111100100110   ;
13'd3139:weight<=16'b0000000000000011   ;
13'd3140:weight<=16'b0000000000010001   ;
13'd3141:weight<=16'b1111111111001000   ;
13'd3142:weight<=16'b1111111111110100   ;
13'd3143:weight<=16'b1111111111100000   ;
13'd3144:weight<=16'b0000000011100100   ;
13'd3145:weight<=16'b0000000001001111   ;
13'd3146:weight<=16'b1111111101101011   ;
13'd3147:weight<=16'b1111111111011010   ;
13'd3148:weight<=16'b0000000001101111   ;
13'd3149:weight<=16'b1111111110001001   ;
13'd3150:weight<=16'b1111111111111011   ;
13'd3151:weight<=16'b1111111101100000   ;
13'd3152:weight<=16'b0000000000111010   ;
13'd3153:weight<=16'b0000000001110011  ;
13'd3154:weight<=16'b0000000011110001   ;
13'd3155:weight<=16'b1111111110101000   ;
13'd3156:weight<=16'b0000000001100000   ;
13'd3157:weight<=16'b1111111110011111   ;
13'd3158:weight<=16'b1111111101001101   ;
13'd3159:weight<=16'b0000000001000000   ;
13'd3160:weight<=16'b0000000000100110   ;
13'd3161:weight<=16'b0000000000011111   ;
13'd3162:weight<=16'b0000000010000101   ;
13'd3163:weight<=16'b1111111111100001   ;
13'd3164:weight<=16'b0000000001011000   ;
13'd3165:weight<=16'b0000000000000011   ;
13'd3166:weight<=16'b1111111110001101   ;
13'd3167:weight<=16'b1111111101001110   ;
13'd3168:weight<=16'b0000000000101000   ;
13'd3169:weight<=16'b1111111111101010   ;
13'd3170:weight<=16'b1111111111101010   ;
13'd3171:weight<=16'b0000000001010010   ;
13'd3172:weight<=16'b0000000001010001   ;
13'd3173:weight<=16'b1111111101011100   ;
13'd3174:weight<=16'b0000000010110100   ;
13'd3175:weight<=16'b0000000010101011   ;
13'd3176:weight<=16'b1111111110110001   ;
13'd3177:weight<=16'b1111111101101000   ;
13'd3178:weight<=16'b1111111111000100   ;
13'd3179:weight<=16'b0000000000000001   ;
13'd3180:weight<=16'b1111111101100100   ;
13'd3181:weight<=16'b0000000000011011   ;
13'd3182:weight<=16'b1111111011110110   ;
13'd3183:weight<=16'b0000000000110001   ;
13'd3184:weight<=16'b1111111110111001   ;
13'd3185:weight<=16'b0000000001001101   ;
13'd3186:weight<=16'b0000000001000000   ;
13'd3187:weight<=16'b0000000100111000   ;
13'd3188:weight<=16'b0000000001011011   ;
13'd3189:weight<=16'b1111111110111101   ;
13'd3190:weight<=16'b0000000000010001   ;
13'd3191:weight<=16'b1111111111001000   ;
13'd3192:weight<=16'b1111111111110100   ;
13'd3193:weight<=16'b1111111111100000   ;
13'd3194:weight<=16'b0000000011100100   ;
13'd3195:weight<=16'b0000000001001111   ;
13'd3196:weight<=16'b1111111101101011   ;
13'd3197:weight<=16'b1111111111011010   ;
13'd3198:weight<=16'b0000000001101111   ;
13'd3199:weight<=16'b1111111110001001   ;
13'd3200:weight<=16'b0000000010001011   ;
13'd3201:weight<=16'b0000000010000010   ;
13'd3202:weight<=16'b0000000001100100   ;
13'd3203:weight<=16'b0000000000010100   ;
13'd3204:weight<=16'b0000000000100001   ;
13'd3205:weight<=16'b0000000000100101   ;
13'd3206:weight<=16'b1111111111111100   ;
13'd3207:weight<=16'b1111111111111010   ;
13'd3208:weight<=16'b1111111110110100   ;
13'd3209:weight<=16'b1111111011101000   ;
13'd3210:weight<=16'b0000000000100110   ;
13'd3211:weight<=16'b0000000000011111   ;
13'd3212:weight<=16'b0000000010000101   ;
13'd3213:weight<=16'b1111111111100001   ;
13'd3214:weight<=16'b0000000001011000   ;
13'd3215:weight<=16'b0000000000000011   ;
13'd3216:weight<=16'b1111111110001101   ;
13'd3217:weight<=16'b1111111101001110   ;
13'd3218:weight<=16'b0000000000101000   ;
13'd3219:weight<=16'b1111111111101010   ;
13'd3220:weight<=16'b0000000001010011   ;
13'd3221:weight<=16'b1111111111100100   ;
13'd3222:weight<=16'b0000000000101001   ;
13'd3223:weight<=16'b0000000011000110   ;
13'd3224:weight<=16'b1111111111100000   ;
13'd3225:weight<=16'b1111111110111101   ;
13'd3226:weight<=16'b0000000000101101   ;
13'd3227:weight<=16'b1111111110011110   ;
13'd3228:weight<=16'b1111111111111001   ;
13'd3229:weight<=16'b1111111110010110   ;
13'd3230:weight<=16'b1111111101100100   ;
13'd3231:weight<=16'b0000000000011011   ;
13'd3232:weight<=16'b1111111011110110   ;
13'd3233:weight<=16'b0000000000110001   ;
13'd3234:weight<=16'b1111111110111001   ;
13'd3235:weight<=16'b0000000001001101   ;
13'd3236:weight<=16'b0000000001000000   ;
13'd3237:weight<=16'b0000000100111000   ;
13'd3238:weight<=16'b0000000001011011   ;
13'd3239:weight<=16'b1111111110111101   ;
13'd3240:weight<=16'b0000000001101110  ;
13'd3241:weight<=16'b0000000010101100   ;
13'd3242:weight<=16'b1111111110111100   ;
13'd3243:weight<=16'b0000000001011010   ;
13'd3244:weight<=16'b1111111101010011   ;
13'd3245:weight<=16'b1111111111101000   ;
13'd3246:weight<=16'b1111111111110101   ;
13'd3247:weight<=16'b1111111101011101   ;
13'd3248:weight<=16'b0000000011001100   ;
13'd3249:weight<=16'b1111111110110010   ;
13'd3250:weight<=16'b0000000010001011   ;
13'd3251:weight<=16'b0000000010000010   ;
13'd3252:weight<=16'b0000000001100100   ;
13'd3253:weight<=16'b0000000000010100   ;
13'd3254:weight<=16'b0000000000100001   ;
13'd3255:weight<=16'b0000000000100101   ;
13'd3256:weight<=16'b1111111111111100   ;
13'd3257:weight<=16'b1111111111111010   ;
13'd3258:weight<=16'b1111111110110100   ;
13'd3259:weight<=16'b1111111011101000   ;
13'd3260:weight<=16'b0000000010010011   ;
13'd3261:weight<=16'b0000000101101011   ;
13'd3262:weight<=16'b1111111110010001   ;
13'd3263:weight<=16'b1111111111000000   ;
13'd3264:weight<=16'b1111111111111100   ;
13'd3265:weight<=16'b1111111110111011   ;
13'd3266:weight<=16'b1111111110100000   ;
13'd3267:weight<=16'b1111111111100010   ;
13'd3268:weight<=16'b0000000001000110   ;
13'd3269:weight<=16'b1111111101000111   ;
13'd3270:weight<=16'b0000000001010011   ;
13'd3271:weight<=16'b1111111111100100   ;
13'd3272:weight<=16'b0000000000101001   ;
13'd3273:weight<=16'b0000000011000110   ;
13'd3274:weight<=16'b1111111111100000   ;
13'd3275:weight<=16'b1111111110111101   ;
13'd3276:weight<=16'b0000000000101101   ;
13'd3277:weight<=16'b1111111110011110   ;
13'd3278:weight<=16'b1111111111111001   ;
13'd3279:weight<=16'b1111111110010110   ;
13'd3280:weight<=16'b0000000001011001   ;
13'd3281:weight<=16'b0000000000010001   ;
13'd3282:weight<=16'b0000000001010100   ;
13'd3283:weight<=16'b1111111111011110   ;
13'd3284:weight<=16'b0000000000101100   ;
13'd3285:weight<=16'b1111111110111110   ;
13'd3286:weight<=16'b0000000000001011   ;
13'd3287:weight<=16'b1111111110110000   ;
13'd3288:weight<=16'b1111111111010111   ;
13'd3289:weight<=16'b0000000000011110   ;
13'd3290:weight<=16'b0000000001101110   ;
13'd3291:weight<=16'b0000000010101100   ;
13'd3292:weight<=16'b1111111110111100   ;
13'd3293:weight<=16'b0000000001011010   ;
13'd3294:weight<=16'b1111111101010011   ;
13'd3295:weight<=16'b1111111111101000   ;
13'd3296:weight<=16'b1111111111110101   ;
13'd3297:weight<=16'b1111111101011101   ;
13'd3298:weight<=16'b0000000011001100   ;
13'd3299:weight<=16'b1111111110110010   ;
13'd3300:weight<=16'b0000000000011111   ;
13'd3301:weight<=16'b0000000001011101   ;
13'd3302:weight<=16'b0000000000011101   ;
13'd3303:weight<=16'b1111111110111100   ;
13'd3304:weight<=16'b1111111110100010   ;
13'd3305:weight<=16'b0000000000000100   ;
13'd3306:weight<=16'b0000000000010100   ;
13'd3307:weight<=16'b1111111111110001   ;
13'd3308:weight<=16'b1111111110001100   ;
13'd3309:weight<=16'b0000000011101111   ;
13'd3310:weight<=16'b0000000010010011   ;
13'd3311:weight<=16'b0000000101101011   ;
13'd3312:weight<=16'b1111111110010001   ;
13'd3313:weight<=16'b1111111111000000   ;
13'd3314:weight<=16'b1111111111111100   ;
13'd3315:weight<=16'b1111111110111011   ;
13'd3316:weight<=16'b1111111110100000   ;
13'd3317:weight<=16'b1111111111100010   ;
13'd3318:weight<=16'b0000000001000110   ;
13'd3319:weight<=16'b1111111101000111   ;
13'd3320:weight<=16'b0000000000110100   ;
13'd3321:weight<=16'b1111111111111100   ;
13'd3322:weight<=16'b0000000100000000   ;
13'd3323:weight<=16'b0000000010001101   ;
13'd3324:weight<=16'b0000000011101101   ;
13'd3325:weight<=16'b0000000011010111   ;
13'd3326:weight<=16'b1111111010000111   ;
13'd3327:weight<=16'b1111111011100001   ;
13'd3328:weight<=16'b0000000000010110   ;
13'd3329:weight<=16'b1111111110001010   ;
13'd3330:weight<=16'b0000000001011001   ;
13'd3331:weight<=16'b0000000000010001   ;
13'd3332:weight<=16'b0000000001010100   ;
13'd3333:weight<=16'b1111111111011110   ;
13'd3334:weight<=16'b0000000000101100   ;
13'd3335:weight<=16'b1111111110111110   ;
13'd3336:weight<=16'b0000000000001011   ;
13'd3337:weight<=16'b1111111110110000   ;
13'd3338:weight<=16'b1111111111010111   ;
13'd3339:weight<=16'b0000000000011110   ;
13'd3340:weight<=16'b0000000001100000   ;
13'd3341:weight<=16'b1111111111010001   ;
13'd3342:weight<=16'b1111111110010011   ;
13'd3343:weight<=16'b0000000001010100   ;
13'd3344:weight<=16'b0000000001001001   ;
13'd3345:weight<=16'b0000000000010101   ;
13'd3346:weight<=16'b1111111101111001   ;
13'd3347:weight<=16'b1111111111101001   ;
13'd3348:weight<=16'b0000000001110101   ;
13'd3349:weight<=16'b1111111110111000   ;
13'd3350:weight<=16'b0000000000011111   ;
13'd3351:weight<=16'b0000000001011101   ;
13'd3352:weight<=16'b0000000000011101   ;
13'd3353:weight<=16'b1111111110111100   ;
13'd3354:weight<=16'b1111111110100010   ;
13'd3355:weight<=16'b0000000000000100   ;
13'd3356:weight<=16'b0000000000010100   ;
13'd3357:weight<=16'b1111111111110001   ;
13'd3358:weight<=16'b1111111110001100   ;
13'd3359:weight<=16'b0000000011101111   ;
13'd3360:weight<=16'b0000000010100100   ;
13'd3361:weight<=16'b0000000001101111   ;
13'd3362:weight<=16'b0000000000101110   ;
13'd3363:weight<=16'b1111111111110111   ;
13'd3364:weight<=16'b1111111111110000   ;
13'd3365:weight<=16'b1111111111011011   ;
13'd3366:weight<=16'b1111111101101010   ;
13'd3367:weight<=16'b1111111101010111   ;
13'd3368:weight<=16'b1111111111110001   ;
13'd3369:weight<=16'b0000000001111010   ;
13'd3370:weight<=16'b0000000000110100   ;
13'd3371:weight<=16'b1111111111111100   ;
13'd3372:weight<=16'b0000000100000000   ;
13'd3373:weight<=16'b0000000010001101   ;
13'd3374:weight<=16'b0000000011101101   ;
13'd3375:weight<=16'b0000000011010111   ;
13'd3376:weight<=16'b1111111010000111   ;
13'd3377:weight<=16'b1111111011100001   ;
13'd3378:weight<=16'b0000000000010110   ;
13'd3379:weight<=16'b1111111110001010   ;
13'd3380:weight<=16'b0000000100110011   ;
13'd3381:weight<=16'b0000000100001011   ;
13'd3382:weight<=16'b1111111101101101   ;
13'd3383:weight<=16'b1111111110110001   ;
13'd3384:weight<=16'b1111111110001001   ;
13'd3385:weight<=16'b0000000001010111   ;
13'd3386:weight<=16'b1111111111000000   ;
13'd3387:weight<=16'b1111111111111000   ;
13'd3388:weight<=16'b1111111111100001   ;
13'd3389:weight<=16'b1111111101010001   ;
13'd3390:weight<=16'b0000000001100000   ;
13'd3391:weight<=16'b1111111111010001   ;
13'd3392:weight<=16'b1111111110010011   ;
13'd3393:weight<=16'b0000000001010100   ;
13'd3394:weight<=16'b0000000001001001   ;
13'd3395:weight<=16'b0000000000010101   ;
13'd3396:weight<=16'b1111111101111001   ;
13'd3397:weight<=16'b1111111111101001   ;
13'd3398:weight<=16'b0000000001110101   ;
13'd3399:weight<=16'b1111111110111000   ;
13'd3400:weight<=16'b0000000001111111   ;
13'd3401:weight<=16'b1111111111000111   ;
13'd3402:weight<=16'b1111111110111110   ;
13'd3403:weight<=16'b0000000011001110   ;
13'd3404:weight<=16'b1111111111001110   ;
13'd3405:weight<=16'b1111111111101100   ;
13'd3406:weight<=16'b0000000000011111   ;
13'd3407:weight<=16'b1111111110100101   ;
13'd3408:weight<=16'b1111111111011101   ;
13'd3409:weight<=16'b1111111111011110   ;
13'd3410:weight<=16'b0000000010100100   ;
13'd3411:weight<=16'b0000000001101111   ;
13'd3412:weight<=16'b0000000000101110   ;
13'd3413:weight<=16'b1111111111110111   ;
13'd3414:weight<=16'b1111111111110000   ;
13'd3415:weight<=16'b1111111111011011   ;
13'd3416:weight<=16'b1111111101101010   ;
13'd3417:weight<=16'b1111111101010111   ;
13'd3418:weight<=16'b1111111111110001   ;
13'd3419:weight<=16'b0000000001111010   ;
13'd3420:weight<=16'b1111111111000111   ;
13'd3421:weight<=16'b0000000001000110   ;
13'd3422:weight<=16'b1111111111001000   ;
13'd3423:weight<=16'b0000000011001101   ;
13'd3424:weight<=16'b0000000000101001   ;
13'd3425:weight<=16'b1111111111101001   ;
13'd3426:weight<=16'b0000000011000100   ;
13'd3427:weight<=16'b0000000001000010   ;
13'd3428:weight<=16'b1111111001001110   ;
13'd3429:weight<=16'b0000000001010110   ;
13'd3430:weight<=16'b0000000100110011   ;
13'd3431:weight<=16'b0000000100001011   ;
13'd3432:weight<=16'b1111111101101101   ;
13'd3433:weight<=16'b1111111110110001   ;
13'd3434:weight<=16'b1111111110001001   ;
13'd3435:weight<=16'b0000000001010111   ;
13'd3436:weight<=16'b1111111111000000   ;
13'd3437:weight<=16'b1111111111111000   ;
13'd3438:weight<=16'b1111111111100001   ;
13'd3439:weight<=16'b1111111101010001   ;
13'd3440:weight<=16'b0000000001000001   ;
13'd3441:weight<=16'b0000000000100100   ;
13'd3442:weight<=16'b0000000000001100   ;
13'd3443:weight<=16'b0000000000011001   ;
13'd3444:weight<=16'b1111111111011111   ;
13'd3445:weight<=16'b0000000001001101   ;
13'd3446:weight<=16'b1111111111010101   ;
13'd3447:weight<=16'b1111111101011010   ;
13'd3448:weight<=16'b0000000001111010   ;
13'd3449:weight<=16'b1111111111010010   ;
13'd3450:weight<=16'b0000000001111111   ;
13'd3451:weight<=16'b1111111111000111   ;
13'd3452:weight<=16'b1111111110111110   ;
13'd3453:weight<=16'b0000000011001110   ;
13'd3454:weight<=16'b1111111111001110   ;
13'd3455:weight<=16'b1111111111101100   ;
13'd3456:weight<=16'b0000000000011111   ;
13'd3457:weight<=16'b1111111110100101   ;
13'd3458:weight<=16'b1111111111011101   ;
13'd3459:weight<=16'b1111111111011110   ;
13'd3460:weight<=16'b0000000001100000   ;
13'd3461:weight<=16'b0000000010000111   ;
13'd3462:weight<=16'b1111111100111110   ;
13'd3463:weight<=16'b0000000011000111   ;
13'd3464:weight<=16'b1111111111111000   ;
13'd3465:weight<=16'b1111111101100100   ;
13'd3466:weight<=16'b0000000000010010   ;
13'd3467:weight<=16'b1111111111001101   ;
13'd3468:weight<=16'b0000000010000101   ;
13'd3469:weight<=16'b1111111110000010   ;
13'd3470:weight<=16'b1111111111000111   ;
13'd3471:weight<=16'b0000000001000110   ;
13'd3472:weight<=16'b1111111111001000   ;
13'd3473:weight<=16'b0000000011001101   ;
13'd3474:weight<=16'b0000000000101001   ;
13'd3475:weight<=16'b1111111111101001   ;
13'd3476:weight<=16'b0000000011000100   ;
13'd3477:weight<=16'b0000000001000010   ;
13'd3478:weight<=16'b1111111001001110   ;
13'd3479:weight<=16'b0000000001010110   ;
13'd3480:weight<=16'b0000000001010101   ;
13'd3481:weight<=16'b0000000010111010   ;
13'd3482:weight<=16'b0000000010110100   ;
13'd3483:weight<=16'b1111111110000000   ;
13'd3484:weight<=16'b0000000000001001   ;
13'd3485:weight<=16'b1111111111100110   ;
13'd3486:weight<=16'b0000000000000100   ;
13'd3487:weight<=16'b0000000001100001   ;
13'd3488:weight<=16'b1111111110000000   ;
13'd3489:weight<=16'b1111111101001001   ;
13'd3490:weight<=16'b0000000001000001   ;
13'd3491:weight<=16'b0000000000100100   ;
13'd3492:weight<=16'b0000000000001100   ;
13'd3493:weight<=16'b0000000000011001   ;
13'd3494:weight<=16'b1111111111011111   ;
13'd3495:weight<=16'b0000000001001101   ;
13'd3496:weight<=16'b1111111111010101   ;
13'd3497:weight<=16'b1111111101011010   ;
13'd3498:weight<=16'b0000000001111010   ;
13'd3499:weight<=16'b1111111111010010   ;
13'd3500:weight<=16'b1111111111011101   ;
13'd3501:weight<=16'b1111111110111001   ;
13'd3502:weight<=16'b0000000001101100   ;
13'd3503:weight<=16'b0000000000110110   ;
13'd3504:weight<=16'b0000000000110010   ;
13'd3505:weight<=16'b1111111111101101   ;
13'd3506:weight<=16'b0000000000110010   ;
13'd3507:weight<=16'b1111111110011000   ;
13'd3508:weight<=16'b1111111111011110   ;
13'd3509:weight<=16'b0000000000110001   ;
13'd3510:weight<=16'b0000000001100000   ;
13'd3511:weight<=16'b0000000010000111   ;
13'd3512:weight<=16'b1111111100111110   ;
13'd3513:weight<=16'b0000000011000111   ;
13'd3514:weight<=16'b1111111111111000   ;
13'd3515:weight<=16'b1111111101100100   ;
13'd3516:weight<=16'b0000000000010010   ;
13'd3517:weight<=16'b1111111111001101   ;
13'd3518:weight<=16'b0000000010000101   ;
13'd3519:weight<=16'b1111111110000010   ;
13'd3520:weight<=16'b1111111111111100   ;
13'd3521:weight<=16'b1111111110101100   ;
13'd3522:weight<=16'b0000000011110010   ;
13'd3523:weight<=16'b0000000000001111   ;
13'd3524:weight<=16'b1111111100110110   ;
13'd3525:weight<=16'b0000000000000011   ;
13'd3526:weight<=16'b0000000000001100  ;
13'd3527:weight<=16'b0000000010011001   ;
13'd3528:weight<=16'b1111111110010000   ;
13'd3529:weight<=16'b0000000001000101   ;
13'd3530:weight<=16'b0000000001010101   ;
13'd3531:weight<=16'b0000000010111010   ;
13'd3532:weight<=16'b0000000010110100   ;
13'd3533:weight<=16'b1111111110000000   ;
13'd3534:weight<=16'b0000000000001001   ;
13'd3535:weight<=16'b1111111111100110   ;
13'd3536:weight<=16'b0000000000000100   ;
13'd3537:weight<=16'b0000000001100001   ;
13'd3538:weight<=16'b1111111110000000   ;
13'd3539:weight<=16'b1111111101001001   ;
13'd3540:weight<=16'b0000000001011011   ;
13'd3541:weight<=16'b0000000001001001   ;
13'd3542:weight<=16'b0000000010101100   ;
13'd3543:weight<=16'b1111111110101011   ;
13'd3544:weight<=16'b1111111110001111   ;
13'd3545:weight<=16'b1111111111000011   ;
13'd3546:weight<=16'b1111111110110111   ;
13'd3547:weight<=16'b0000000001101011   ;
13'd3548:weight<=16'b1111111110000101   ;
13'd3549:weight<=16'b0000000000101011   ;
13'd3550:weight<=16'b1111111111011101   ;
13'd3551:weight<=16'b1111111110111001   ;
13'd3552:weight<=16'b0000000001101100   ;
13'd3553:weight<=16'b0000000000110110   ;
13'd3554:weight<=16'b0000000000110010   ;
13'd3555:weight<=16'b1111111111101101   ;
13'd3556:weight<=16'b0000000000110010   ;
13'd3557:weight<=16'b1111111110011000   ;
13'd3558:weight<=16'b1111111111011110   ;
13'd3559:weight<=16'b0000000000110001   ;
13'd3560:weight<=16'b0000000001001001   ;
13'd3561:weight<=16'b0000000100000001   ;
13'd3562:weight<=16'b1111111100000011   ;
13'd3563:weight<=16'b0000000110110100   ;
13'd3564:weight<=16'b1111111000110101   ;
13'd3565:weight<=16'b0000000011000100   ;
13'd3566:weight<=16'b1111110110100110   ;
13'd3567:weight<=16'b0000000101011101   ;
13'd3568:weight<=16'b0000000100100100   ;
13'd3569:weight<=16'b1111111001110011   ;
13'd3570:weight<=16'b1111111111111100   ;
13'd3571:weight<=16'b1111111110101100   ;
13'd3572:weight<=16'b0000000011110010   ;
13'd3573:weight<=16'b0000000000001111   ;
13'd3574:weight<=16'b1111111100110110   ;
13'd3575:weight<=16'b0000000000000011   ;
13'd3576:weight<=16'b0000000000001100   ;
13'd3577:weight<=16'b0000000010011001   ;
13'd3578:weight<=16'b1111111110010000   ;
13'd3579:weight<=16'b0000000001000101   ;
13'd3580:weight<=16'b0000000010110010   ;
13'd3581:weight<=16'b0000000010001101   ;
13'd3582:weight<=16'b1111111010010010   ;
13'd3583:weight<=16'b0000000010100011   ;
13'd3584:weight<=16'b1111111101111100   ;
13'd3585:weight<=16'b0000000110001011   ;
13'd3586:weight<=16'b0000000010100010   ;
13'd3587:weight<=16'b1111111100001000   ;
13'd3588:weight<=16'b0000000000111010   ;
13'd3589:weight<=16'b1111111100011110   ;
13'd3590:weight<=16'b0000000001011011   ;
13'd3591:weight<=16'b0000000001001001   ;
13'd3592:weight<=16'b0000000010101100   ;
13'd3593:weight<=16'b1111111110101011   ;
13'd3594:weight<=16'b1111111110001111   ;
13'd3595:weight<=16'b1111111111000011   ;
13'd3596:weight<=16'b1111111110110111   ;
13'd3597:weight<=16'b0000000001101011   ;
13'd3598:weight<=16'b1111111110000101   ;
13'd3599:weight<=16'b0000000000101011   ;
13'd3600:weight<=16'b1111111110011100   ;
13'd3601:weight<=16'b1111111111000010   ;
13'd3602:weight<=16'b1111111111010111   ;
13'd3603:weight<=16'b0000000001000011   ;
13'd3604:weight<=16'b0000000001100100   ;
13'd3605:weight<=16'b0000000010100110   ;
13'd3606:weight<=16'b1111111111100100   ;
13'd3607:weight<=16'b1111111110101100   ;
13'd3608:weight<=16'b1111111111111010   ;
13'd3609:weight<=16'b0000000000011100   ;
13'd3610:weight<=16'b0000000001001001   ;
13'd3611:weight<=16'b0000000100000001   ;
13'd3612:weight<=16'b1111111100000011   ;
13'd3613:weight<=16'b0000000110110100   ;
13'd3614:weight<=16'b1111111000110101   ;
13'd3615:weight<=16'b0000000011000100   ;
13'd3616:weight<=16'b1111110110100110   ;
13'd3617:weight<=16'b0000000101011101   ;
13'd3618:weight<=16'b0000000100100100   ;
13'd3619:weight<=16'b1111111001110011   ;
13'd3620:weight<=16'b0000000001001001   ;
13'd3621:weight<=16'b1111111111111010   ;
13'd3622:weight<=16'b1111111111011111   ;
13'd3623:weight<=16'b0000000000000010   ;
13'd3624:weight<=16'b1111111111110011   ;
13'd3625:weight<=16'b1111111110101111   ;
13'd3626:weight<=16'b0000000000111100   ;
13'd3627:weight<=16'b1111111111110101   ;
13'd3628:weight<=16'b0000000001010010   ;
13'd3629:weight<=16'b1111111110100001   ;
13'd3630:weight<=16'b0000000010110010   ;
13'd3631:weight<=16'b0000000010001101   ;
13'd3632:weight<=16'b1111111010010010   ;
13'd3633:weight<=16'b0000000010100011   ;
13'd3634:weight<=16'b1111111101111100   ;
13'd3635:weight<=16'b0000000110001011   ;
13'd3636:weight<=16'b0000000010100010   ;
13'd3637:weight<=16'b1111111100001000   ;
13'd3638:weight<=16'b0000000000111010   ;
13'd3639:weight<=16'b1111111100011110   ;
13'd3640:weight<=16'b0000000001010101   ;
13'd3641:weight<=16'b1111111111111011   ;
13'd3642:weight<=16'b1111111101011011   ;
13'd3643:weight<=16'b1111111111111011   ;
13'd3644:weight<=16'b1111111110011011   ;
13'd3645:weight<=16'b0000000000010001   ;
13'd3646:weight<=16'b0000000001000100   ;
13'd3647:weight<=16'b0000000000101000   ;
13'd3648:weight<=16'b0000000000110001   ;
13'd3649:weight<=16'b1111111111111011   ;
13'd3650:weight<=16'b1111111110011100   ;
13'd3651:weight<=16'b1111111111000010   ;
13'd3652:weight<=16'b1111111111010111   ;
13'd3653:weight<=16'b0000000001000011   ;
13'd3654:weight<=16'b0000000001100100   ;
13'd3655:weight<=16'b0000000010100110   ;
13'd3656:weight<=16'b1111111111100100   ;
13'd3657:weight<=16'b1111111110101100   ;
13'd3658:weight<=16'b1111111111111010   ;
13'd3659:weight<=16'b0000000000011100   ;
13'd3660:weight<=16'b0000000000111110   ;
13'd3661:weight<=16'b0000000010001110   ;
13'd3662:weight<=16'b1111111110110001   ;
13'd3663:weight<=16'b0000000010001101   ;
13'd3664:weight<=16'b1111111111111000   ;
13'd3665:weight<=16'b0000000000011111   ;
13'd3666:weight<=16'b1111111101110010   ;
13'd3667:weight<=16'b1111111110100001   ;
13'd3668:weight<=16'b1111111111010101   ;
13'd3669:weight<=16'b1111111111111010   ;
13'd3670:weight<=16'b0000000001001001   ;
13'd3671:weight<=16'b1111111111111010   ;
13'd3672:weight<=16'b1111111111011111   ;
13'd3673:weight<=16'b0000000000000010   ;
13'd3674:weight<=16'b1111111111110011   ;
13'd3675:weight<=16'b1111111110101111   ;
13'd3676:weight<=16'b0000000000111100   ;
13'd3677:weight<=16'b1111111111110101   ;
13'd3678:weight<=16'b0000000001010010   ;
13'd3679:weight<=16'b1111111110100001   ;
13'd3680:weight<=16'b0000000000000000   ;
13'd3681:weight<=16'b0000000000101111   ;
13'd3682:weight<=16'b0000000000010011   ;
13'd3683:weight<=16'b1111111101110010   ;
13'd3684:weight<=16'b0000000000011110   ;
13'd3685:weight<=16'b0000000010100001   ;
13'd3686:weight<=16'b0000000000011001   ;
13'd3687:weight<=16'b1111111111111011   ;
13'd3688:weight<=16'b1111111101010010   ;
13'd3689:weight<=16'b0000000001101001   ;
13'd3690:weight<=16'b0000000001010101   ;
13'd3691:weight<=16'b1111111111111011   ;
13'd3692:weight<=16'b1111111101011011   ;
13'd3693:weight<=16'b1111111111111011   ;
13'd3694:weight<=16'b1111111110011011  ;
13'd3695:weight<=16'b0000000000010001   ;
13'd3696:weight<=16'b0000000001000100   ;
13'd3697:weight<=16'b0000000000101000   ;
13'd3698:weight<=16'b0000000000110001   ;
13'd3699:weight<=16'b1111111111111011   ;
13'd3700:weight<=16'b0000000001101010   ;
13'd3701:weight<=16'b0000000000101100   ;
13'd3702:weight<=16'b0000000001010000   ;
13'd3703:weight<=16'b0000000000010101   ;
13'd3704:weight<=16'b1111111111010100   ;
13'd3705:weight<=16'b1111111110100101   ;
13'd3706:weight<=16'b0000000000010100   ;
13'd3707:weight<=16'b1111111111001111   ;
13'd3708:weight<=16'b1111111110101100   ;
13'd3709:weight<=16'b0000000000010000   ;
13'd3710:weight<=16'b0000000000111110   ;
13'd3711:weight<=16'b0000000010001110   ;
13'd3712:weight<=16'b1111111110110001   ;
13'd3713:weight<=16'b0000000010001101   ;
13'd3714:weight<=16'b1111111111111000   ;
13'd3715:weight<=16'b0000000000011111   ;
13'd3716:weight<=16'b1111111101110010   ;
13'd3717:weight<=16'b1111111110100001   ;
13'd3718:weight<=16'b1111111111010101   ;
13'd3719:weight<=16'b1111111111111010   ;
13'd3720:weight<=16'b1111111110111110   ;
13'd3721:weight<=16'b0000000000000100   ;
13'd3722:weight<=16'b1111111110100001   ;
13'd3723:weight<=16'b0000000000101110   ;
13'd3724:weight<=16'b1111111111100110   ;
13'd3725:weight<=16'b0000000010001001   ;
13'd3726:weight<=16'b0000000001001100   ;
13'd3727:weight<=16'b1111111111101101   ;
13'd3728:weight<=16'b0000000000111110   ;
13'd3729:weight<=16'b1111111110101000   ;
13'd3730:weight<=16'b0000000000000000   ;
13'd3731:weight<=16'b0000000000101111   ;
13'd3732:weight<=16'b0000000000010011   ;
13'd3733:weight<=16'b1111111101110010   ;
13'd3734:weight<=16'b0000000000011110   ;
13'd3735:weight<=16'b0000000010100001   ;
13'd3736:weight<=16'b0000000000011001   ;
13'd3737:weight<=16'b1111111111111011   ;
13'd3738:weight<=16'b1111111101010010   ;
13'd3739:weight<=16'b0000000001101001   ;
13'd3740:weight<=16'b0000000000000001   ;
13'd3741:weight<=16'b1111111110110001   ;
13'd3742:weight<=16'b1111111111110110   ;
13'd3743:weight<=16'b1111111111101011   ;
13'd3744:weight<=16'b0000000000011001   ;
13'd3745:weight<=16'b1111111111011110   ;
13'd3746:weight<=16'b1111111111101110   ;
13'd3747:weight<=16'b0000000001001101   ;
13'd3748:weight<=16'b0000000000011000   ;
13'd3749:weight<=16'b0000000000110001   ;
13'd3750:weight<=16'b0000000001101010   ;
13'd3751:weight<=16'b0000000000101100   ;
13'd3752:weight<=16'b0000000001010000   ;
13'd3753:weight<=16'b0000000000010101   ;
13'd3754:weight<=16'b1111111111010100   ;
13'd3755:weight<=16'b1111111110100101   ;
13'd3756:weight<=16'b0000000000010100   ;
13'd3757:weight<=16'b1111111111001111   ;
13'd3758:weight<=16'b1111111110101100   ;
13'd3759:weight<=16'b0000000000010000   ;
13'd3760:weight<=16'b1111111101110111   ;
13'd3761:weight<=16'b1111111111110011   ;
13'd3762:weight<=16'b1111111111000001   ;
13'd3763:weight<=16'b0000000000010100   ;
13'd3764:weight<=16'b0000000000101000   ;
13'd3765:weight<=16'b0000000000010100   ;
13'd3766:weight<=16'b0000000001011010   ;
13'd3767:weight<=16'b1111111111011111   ;
13'd3768:weight<=16'b0000000001111101   ;
13'd3769:weight<=16'b1111111111010010   ;
13'd3770:weight<=16'b1111111110111110   ;
13'd3771:weight<=16'b0000000000000100   ;
13'd3772:weight<=16'b1111111110100001   ;
13'd3773:weight<=16'b0000000000101110   ;
13'd3774:weight<=16'b1111111111100110   ;
13'd3775:weight<=16'b0000000010001001   ;
13'd3776:weight<=16'b0000000001001100   ;
13'd3777:weight<=16'b1111111111101101   ;
13'd3778:weight<=16'b0000000000111110   ;
13'd3779:weight<=16'b1111111110101000   ;
13'd3780:weight<=16'b1111111101000001   ;
13'd3781:weight<=16'b0000000010010011   ;
13'd3782:weight<=16'b1111111010011010   ;
13'd3783:weight<=16'b1111111111110101   ;
13'd3784:weight<=16'b0000000111011010   ;
13'd3785:weight<=16'b0000000000110010   ;
13'd3786:weight<=16'b1111111110110101   ;
13'd3787:weight<=16'b1111111111110111   ;
13'd3788:weight<=16'b1111111111001001   ;
13'd3789:weight<=16'b0000000010101000   ;
13'd3790:weight<=16'b0000000000000001   ;
13'd3791:weight<=16'b1111111110110001   ;
13'd3792:weight<=16'b1111111111110110   ;
13'd3793:weight<=16'b1111111111101011   ;
13'd3794:weight<=16'b0000000000011001   ;
13'd3795:weight<=16'b1111111111011110   ;
13'd3796:weight<=16'b1111111111101110   ;
13'd3797:weight<=16'b0000000001001101   ;
13'd3798:weight<=16'b0000000000011000   ;
13'd3799:weight<=16'b0000000000110001   ;
13'd3800:weight<=16'b1111111111000110   ;
13'd3801:weight<=16'b0000000011000010   ;
13'd3802:weight<=16'b1111111101101010   ;
13'd3803:weight<=16'b0000000111101010   ;
13'd3804:weight<=16'b0000000000000001   ;
13'd3805:weight<=16'b1111111100001000   ;
13'd3806:weight<=16'b0000000011011100   ;
13'd3807:weight<=16'b1111111110101001   ;
13'd3808:weight<=16'b1111111010110110   ;
13'd3809:weight<=16'b0000000000001010   ;
13'd3810:weight<=16'b1111111101110111   ;
13'd3811:weight<=16'b1111111111110011   ;
13'd3812:weight<=16'b1111111111000001   ;
13'd3813:weight<=16'b0000000000010100   ;
13'd3814:weight<=16'b0000000000101000   ;
13'd3815:weight<=16'b0000000000010100   ;
13'd3816:weight<=16'b0000000001011010   ;
13'd3817:weight<=16'b1111111111011111   ;
13'd3818:weight<=16'b0000000001111101   ;
13'd3819:weight<=16'b1111111111010010   ;
13'd3820:weight<=16'b0000000001110010   ;
13'd3821:weight<=16'b0000000010101001   ;
13'd3822:weight<=16'b1111111110010110   ;
13'd3823:weight<=16'b1111111111100001   ;
13'd3824:weight<=16'b1111111110100111   ;
13'd3825:weight<=16'b1111111101100111   ;
13'd3826:weight<=16'b1111111101101110   ;
13'd3827:weight<=16'b0000000110011100   ;
13'd3828:weight<=16'b1111111100110110   ;
13'd3829:weight<=16'b0000000001010001   ;
13'd3830:weight<=16'b1111111101000001   ;
13'd3831:weight<=16'b0000000010010011   ;
13'd3832:weight<=16'b1111111010011010   ;
13'd3833:weight<=16'b1111111111110101   ;
13'd3834:weight<=16'b0000000111011010   ;
13'd3835:weight<=16'b0000000000110010   ;
13'd3836:weight<=16'b1111111110110101   ;
13'd3837:weight<=16'b1111111111110111   ;
13'd3838:weight<=16'b1111111111001001   ;
13'd3839:weight<=16'b0000000010101000   ;
13'd3840:weight<=16'b1111111010101011   ;
13'd3841:weight<=16'b1111111100101110   ;
13'd3842:weight<=16'b0000000111110001   ;
13'd3843:weight<=16'b1111111101111111   ;
13'd3844:weight<=16'b1111111110000100   ;
13'd3845:weight<=16'b0000001000010001   ;
13'd3846:weight<=16'b1111111110001101   ;
13'd3847:weight<=16'b0000000100010111   ;
13'd3848:weight<=16'b1111111100101101   ;
13'd3849:weight<=16'b1111111110111110   ;
13'd3850:weight<=16'b1111111111000110   ;
13'd3851:weight<=16'b0000000011000010   ;
13'd3852:weight<=16'b1111111101101010   ;
13'd3853:weight<=16'b0000000111101010   ;
13'd3854:weight<=16'b0000000000000001   ;
13'd3855:weight<=16'b1111111100001000   ;
13'd3856:weight<=16'b0000000011011100   ;
13'd3857:weight<=16'b1111111110101001   ;
13'd3858:weight<=16'b1111111010110110   ;
13'd3859:weight<=16'b0000000000001010   ;
13'd3860:weight<=16'b1111111100010001   ;
13'd3861:weight<=16'b0000000001001001   ;
13'd3862:weight<=16'b1111111111001101   ;
13'd3863:weight<=16'b0000000001001100   ;
13'd3864:weight<=16'b0000000001110101   ;
13'd3865:weight<=16'b0000000001001101   ;
13'd3866:weight<=16'b0000000101001111   ;
13'd3867:weight<=16'b1111111111001000   ;
13'd3868:weight<=16'b1111111011010011   ;
13'd3869:weight<=16'b0000000000111011   ;
13'd3870:weight<=16'b0000000001110010   ;
13'd3871:weight<=16'b0000000010101001   ;
13'd3872:weight<=16'b1111111110010110   ;
13'd3873:weight<=16'b1111111111100001   ;
13'd3874:weight<=16'b1111111110100111   ;
13'd3875:weight<=16'b1111111101100111   ;
13'd3876:weight<=16'b1111111101101110   ;
13'd3877:weight<=16'b0000000110011100   ;
13'd3878:weight<=16'b1111111100110110   ;
13'd3879:weight<=16'b0000000001010001   ;
13'd3880:weight<=16'b0000000000010101   ;
13'd3881:weight<=16'b1111111111001100   ;
13'd3882:weight<=16'b0000000000010110   ;
13'd3883:weight<=16'b0000000000101000   ;
13'd3884:weight<=16'b1111111111011000   ;
13'd3885:weight<=16'b1111111111110001   ;
13'd3886:weight<=16'b0000000000110110   ;
13'd3887:weight<=16'b0000000010000111   ;
13'd3888:weight<=16'b1111111100010101   ;
13'd3889:weight<=16'b0000000001100011   ;
13'd3890:weight<=16'b1111111010101011   ;
13'd3891:weight<=16'b1111111100101110   ;
13'd3892:weight<=16'b0000000111110001   ;
13'd3893:weight<=16'b1111111101111111   ;
13'd3894:weight<=16'b1111111110000100   ;
13'd3895:weight<=16'b0000001000010001   ;
13'd3896:weight<=16'b1111111110001101   ;
13'd3897:weight<=16'b0000000100010111   ;
13'd3898:weight<=16'b1111111100101101   ;
13'd3899:weight<=16'b1111111110111110   ;
13'd3900:weight<=16'b1111111110011011   ;
13'd3901:weight<=16'b1111111110111000   ;
13'd3902:weight<=16'b0000000001001100   ;
13'd3903:weight<=16'b1111111111101101   ;
13'd3904:weight<=16'b0000000100111000   ;
13'd3905:weight<=16'b1111111101111101   ;
13'd3906:weight<=16'b1111111111111010   ;
13'd3907:weight<=16'b1111111110111100   ;
13'd3908:weight<=16'b1111111100101111   ;
13'd3909:weight<=16'b0000000011110101   ;
13'd3910:weight<=16'b1111111100010001   ;
13'd3911:weight<=16'b0000000001001001   ;
13'd3912:weight<=16'b1111111111001101   ;
13'd3913:weight<=16'b0000000001001100   ;
13'd3914:weight<=16'b0000000001110101   ;
13'd3915:weight<=16'b0000000001001101   ;
13'd3916:weight<=16'b0000000101001111   ;
13'd3917:weight<=16'b1111111111001000   ;
13'd3918:weight<=16'b1111111011010011   ;
13'd3919:weight<=16'b0000000000111011   ;
13'd3920:weight<=16'b1111111111100101   ;
13'd3921:weight<=16'b1111111111011010   ;
13'd3922:weight<=16'b1111111110011000   ;
13'd3923:weight<=16'b0000000000010000   ;
13'd3924:weight<=16'b0000000000101000   ;
13'd3925:weight<=16'b0000000000001010   ;
13'd3926:weight<=16'b1111111110010011   ;
13'd3927:weight<=16'b1111111110000100   ;
13'd3928:weight<=16'b0000000000101100   ;
13'd3929:weight<=16'b0000000100000010   ;
13'd3930:weight<=16'b0000000000010101   ;
13'd3931:weight<=16'b1111111111001100   ;
13'd3932:weight<=16'b0000000000010110   ;
13'd3933:weight<=16'b0000000000101000   ;
13'd3934:weight<=16'b1111111111011000   ;
13'd3935:weight<=16'b1111111111110001   ;
13'd3936:weight<=16'b0000000000110110   ;
13'd3937:weight<=16'b0000000010000111   ;
13'd3938:weight<=16'b1111111100010101   ;
13'd3939:weight<=16'b0000000001100011   ;
13'd3940:weight<=16'b0000000000101011   ;
13'd3941:weight<=16'b0000000011001001   ;
13'd3942:weight<=16'b1111111111000000   ;
13'd3943:weight<=16'b0000000000000011   ;
13'd3944:weight<=16'b1111111110100100   ;
13'd3945:weight<=16'b1111111110001011   ;
13'd3946:weight<=16'b1111111110000111   ;
13'd3947:weight<=16'b1111111110110011   ;
13'd3948:weight<=16'b0000000001001011   ;
13'd3949:weight<=16'b0000000010101011   ;
13'd3950:weight<=16'b1111111110011011   ;
13'd3951:weight<=16'b1111111110111000   ;
13'd3952:weight<=16'b0000000001001100   ;
13'd3953:weight<=16'b1111111111101101   ;
13'd3954:weight<=16'b0000000100111000   ;
13'd3955:weight<=16'b1111111101111101   ;
13'd3956:weight<=16'b1111111111111010   ;
13'd3957:weight<=16'b1111111110111100   ;
13'd3958:weight<=16'b1111111100101111   ;
13'd3959:weight<=16'b0000000011110101   ;
13'd3960:weight<=16'b1111111110111111   ;
13'd3961:weight<=16'b1111111101000101   ;
13'd3962:weight<=16'b0000000010001101   ;
13'd3963:weight<=16'b0000000010100011   ;
13'd3964:weight<=16'b0000000001101100   ;
13'd3965:weight<=16'b1111111110000101   ;
13'd3966:weight<=16'b0000000010010100   ;
13'd3967:weight<=16'b0000000001011110   ;
13'd3968:weight<=16'b1111111011001001   ;
13'd3969:weight<=16'b0000000011110110   ;
13'd3970:weight<=16'b1111111111100101   ;
13'd3971:weight<=16'b1111111111011010   ;
13'd3972:weight<=16'b1111111110011000   ;
13'd3973:weight<=16'b0000000000010000   ;
13'd3974:weight<=16'b0000000000101000   ;
13'd3975:weight<=16'b0000000000001010   ;
13'd3976:weight<=16'b1111111110010011   ;
13'd3977:weight<=16'b1111111110000100   ;
13'd3978:weight<=16'b0000000000101100   ;
13'd3979:weight<=16'b0000000100000010   ;
13'd3980:weight<=16'b0000000001010010   ;
13'd3981:weight<=16'b0000000010101011   ;
13'd3982:weight<=16'b1111111111111010   ;
13'd3983:weight<=16'b1111111101100111   ;
13'd3984:weight<=16'b1111111100011000   ;
13'd3985:weight<=16'b0000000011101101   ;
13'd3986:weight<=16'b1111111110110101   ;
13'd3987:weight<=16'b1111111110001010   ;
13'd3988:weight<=16'b0000000001010111   ;
13'd3989:weight<=16'b0000000010010111   ;
13'd3990:weight<=16'b0000000000101011   ;
13'd3991:weight<=16'b0000000011001001   ;
13'd3992:weight<=16'b1111111111000000   ;
13'd3993:weight<=16'b0000000000000011   ;
13'd3994:weight<=16'b1111111110100100   ;
13'd3995:weight<=16'b1111111110001011   ;
13'd3996:weight<=16'b1111111110000111   ;
13'd3997:weight<=16'b1111111110110011   ;
13'd3998:weight<=16'b0000000001001011   ;
13'd3999:weight<=16'b0000000010101011   ;
13'd4000:weight<=16'b0000000110001000   ;
13'd4001:weight<=16'b1111111110011011   ;
13'd4002:weight<=16'b0000000011001111   ;
13'd4003:weight<=16'b1111111101011011   ;
13'd4004:weight<=16'b1111111110101001   ;
13'd4005:weight<=16'b0000000001111101   ;
13'd4006:weight<=16'b1111111101111011   ;
13'd4007:weight<=16'b0000000000110010   ;
13'd4008:weight<=16'b1111111010001010   ;
13'd4009:weight<=16'b0000000010000010   ;
13'd4010:weight<=16'b1111111110111111   ;
13'd4011:weight<=16'b1111111101000101   ;
13'd4012:weight<=16'b0000000010001101   ;
13'd4013:weight<=16'b0000000010100011   ;
13'd4014:weight<=16'b0000000001101100   ;
13'd4015:weight<=16'b1111111110000101   ;
13'd4016:weight<=16'b0000000010010100   ;
13'd4017:weight<=16'b0000000001011110   ;
13'd4018:weight<=16'b1111111011001001   ;
13'd4019:weight<=16'b0000000011110110   ;
13'd4020:weight<=16'b1111111111000010   ;
13'd4021:weight<=16'b1111111110101010   ;
13'd4022:weight<=16'b0000000001100100   ;
13'd4023:weight<=16'b1111111100111101   ;
13'd4024:weight<=16'b0000000001010011   ;
13'd4025:weight<=16'b0000000001010011   ;
13'd4026:weight<=16'b1111111111111100   ;
13'd4027:weight<=16'b1111111101111001   ;
13'd4028:weight<=16'b0000000010111010   ;
13'd4029:weight<=16'b0000000000011101   ;
13'd4030:weight<=16'b0000000001010010   ;
13'd4031:weight<=16'b0000000010101011   ;
13'd4032:weight<=16'b1111111111111010   ;
13'd4033:weight<=16'b1111111101100111   ;
13'd4034:weight<=16'b1111111100011000   ;
13'd4035:weight<=16'b0000000011101101   ;
13'd4036:weight<=16'b1111111110110101   ;
13'd4037:weight<=16'b1111111110001010   ;
13'd4038:weight<=16'b0000000001010111   ;
13'd4039:weight<=16'b0000000010010111   ;
13'd4040:weight<=16'b0000000000111010   ;
13'd4041:weight<=16'b1111111111011100   ;
13'd4042:weight<=16'b1111111111110010   ;
13'd4043:weight<=16'b1111111111101101   ;
13'd4044:weight<=16'b1111111100110100   ;
13'd4045:weight<=16'b0000000001101011   ;
13'd4046:weight<=16'b1111111111101001   ;
13'd4047:weight<=16'b0000000000111000   ;
13'd4048:weight<=16'b0000000000100000   ;
13'd4049:weight<=16'b0000000000101010   ;
13'd4050:weight<=16'b0000000110001000   ;
13'd4051:weight<=16'b1111111110011011   ;
13'd4052:weight<=16'b0000000011001111   ;
13'd4053:weight<=16'b1111111101011011   ;
13'd4054:weight<=16'b1111111110101001   ;
13'd4055:weight<=16'b0000000001111101   ;
13'd4056:weight<=16'b1111111101111011   ;
13'd4057:weight<=16'b0000000000110010   ;
13'd4058:weight<=16'b1111111010001010   ;
13'd4059:weight<=16'b0000000010000010   ;
13'd4060:weight<=16'b0000000001001111   ;
13'd4061:weight<=16'b1111110100101101   ;
13'd4062:weight<=16'b0000000100000011   ;
13'd4063:weight<=16'b1111111000110101   ;
13'd4064:weight<=16'b0000000000110001   ;
13'd4065:weight<=16'b1111111100011101   ;
13'd4066:weight<=16'b0000001001011001   ;
13'd4067:weight<=16'b1111111100100001   ;
13'd4068:weight<=16'b0000000001010100   ;
13'd4069:weight<=16'b0000000101001101   ;
13'd4070:weight<=16'b1111111111000010   ;
13'd4071:weight<=16'b1111111110101010   ;
13'd4072:weight<=16'b0000000001100100   ;
13'd4073:weight<=16'b1111111100111101   ;
13'd4074:weight<=16'b0000000001010011   ;
13'd4075:weight<=16'b0000000001010011   ;
13'd4076:weight<=16'b1111111111111100   ;
13'd4077:weight<=16'b1111111101111001   ;
13'd4078:weight<=16'b0000000010111010   ;
13'd4079:weight<=16'b0000000000011101   ;
13'd4080:weight<=16'b1111111101111101   ;
13'd4081:weight<=16'b0000000001011010   ;
13'd4082:weight<=16'b1111111110011111   ;
13'd4083:weight<=16'b1111111111110000   ;
13'd4084:weight<=16'b1111111110101001   ;
13'd4085:weight<=16'b0000000000001000   ;
13'd4086:weight<=16'b0000000010101111   ;
13'd4087:weight<=16'b1111111111100100   ;
13'd4088:weight<=16'b0000000001111000   ;
13'd4089:weight<=16'b1111111111001000   ;
13'd4090:weight<=16'b0000000000111010   ;
13'd4091:weight<=16'b1111111111011100   ;
13'd4092:weight<=16'b1111111111110010   ;
13'd4093:weight<=16'b1111111111101101   ;
13'd4094:weight<=16'b1111111100110100   ;
13'd4095:weight<=16'b0000000001101011   ;
13'd4096:weight<=16'b1111111111101001   ;
13'd4097:weight<=16'b0000000000111000   ;
13'd4098:weight<=16'b0000000000100000   ;
13'd4099:weight<=16'b0000000000101010   ;
13'd4100:weight<=16'b1111111110101011   ;
13'd4101:weight<=16'b0000000000011000   ;
13'd4102:weight<=16'b1111111110101110   ;
13'd4103:weight<=16'b0000000000110111   ;
13'd4104:weight<=16'b1111111110000001   ;
13'd4105:weight<=16'b1111111111010100   ;
13'd4106:weight<=16'b0000000011100111   ;
13'd4107:weight<=16'b0000000101000011   ;
13'd4108:weight<=16'b0000000000000101   ;
13'd4109:weight<=16'b1111111101100110   ;
13'd4110:weight<=16'b0000000001001111   ;
13'd4111:weight<=16'b1111110100101101   ;
13'd4112:weight<=16'b0000000100000011   ;
13'd4113:weight<=16'b1111111000110101   ;
13'd4114:weight<=16'b0000000000110001   ;
13'd4115:weight<=16'b1111111100011101   ;
13'd4116:weight<=16'b0000001001011001   ;
13'd4117:weight<=16'b1111111100100001   ;
13'd4118:weight<=16'b0000000001010100   ;
13'd4119:weight<=16'b0000000101001101   ;
13'd4120:weight<=16'b0000000000100001   ;
13'd4121:weight<=16'b1111111101010101   ;
13'd4122:weight<=16'b1111111111110100   ;
13'd4123:weight<=16'b0000000011001001   ;
13'd4124:weight<=16'b0000000000001001   ;
13'd4125:weight<=16'b1111111101001011   ;
13'd4126:weight<=16'b0000000010011101   ;
13'd4127:weight<=16'b0000000000011101   ;
13'd4128:weight<=16'b0000000010100111   ;
13'd4129:weight<=16'b1111111101011001   ;
13'd4130:weight<=16'b1111111101111101   ;
13'd4131:weight<=16'b0000000001011010   ;
13'd4132:weight<=16'b1111111110011111   ;
13'd4133:weight<=16'b1111111111110000   ;
13'd4134:weight<=16'b1111111110101001   ;
13'd4135:weight<=16'b0000000000001000   ;
13'd4136:weight<=16'b0000000010101111   ;
13'd4137:weight<=16'b1111111111100100   ;
13'd4138:weight<=16'b0000000001111000   ;
13'd4139:weight<=16'b1111111111001000   ;
13'd4140:weight<=16'b0000000000101111   ;
13'd4141:weight<=16'b1111111101100110   ;
13'd4142:weight<=16'b1111111110001110   ;
13'd4143:weight<=16'b0000000011010001   ;
13'd4144:weight<=16'b1111111111001010  ;
13'd4145:weight<=16'b1111111110011011   ;
13'd4146:weight<=16'b1111111110011110   ;
13'd4147:weight<=16'b0000000000000100   ;
13'd4148:weight<=16'b0000000010111010   ;
13'd4149:weight<=16'b0000000001010001   ;
13'd4150:weight<=16'b1111111110101011   ;
13'd4151:weight<=16'b0000000000011000   ;
13'd4152:weight<=16'b1111111110101110   ;
13'd4153:weight<=16'b0000000000110111   ;
13'd4154:weight<=16'b1111111110000001   ;
13'd4155:weight<=16'b1111111111010100   ;
13'd4156:weight<=16'b0000000011100111   ;
13'd4157:weight<=16'b0000000101000011   ;
13'd4158:weight<=16'b0000000000000101   ;
13'd4159:weight<=16'b1111111101100110   ;
13'd4160:weight<=16'b0000000000110101   ;
13'd4161:weight<=16'b1111111110010101   ;
13'd4162:weight<=16'b0000000000100110   ;
13'd4163:weight<=16'b1111111111010000   ;
13'd4164:weight<=16'b0000000001111011   ;
13'd4165:weight<=16'b1111111111110001   ;
13'd4166:weight<=16'b1111111100001011   ;
13'd4167:weight<=16'b0000000010000110   ;
13'd4168:weight<=16'b0000000010100010   ;
13'd4169:weight<=16'b1111111111101000   ;
13'd4170:weight<=16'b0000000000100001   ;
13'd4171:weight<=16'b1111111101010101   ;
13'd4172:weight<=16'b1111111111110100   ;
13'd4173:weight<=16'b0000000011001001   ;
13'd4174:weight<=16'b0000000000001001   ;
13'd4175:weight<=16'b1111111101001011   ;
13'd4176:weight<=16'b0000000010011101   ;
13'd4177:weight<=16'b0000000000011101   ;
13'd4178:weight<=16'b0000000010100111   ;
13'd4179:weight<=16'b1111111101011001   ;
13'd4180:weight<=16'b0000000000000011   ;
13'd4181:weight<=16'b0000000000001011   ;
13'd4182:weight<=16'b1111111110100100   ;
13'd4183:weight<=16'b1111111101011100   ;
13'd4184:weight<=16'b0000000000111100   ;
13'd4185:weight<=16'b0000000000010000   ;
13'd4186:weight<=16'b0000000001101000   ;
13'd4187:weight<=16'b0000000001000010   ;
13'd4188:weight<=16'b0000000010011001   ;
13'd4189:weight<=16'b1111111101100011   ;
13'd4190:weight<=16'b0000000000101111   ;
13'd4191:weight<=16'b1111111101100110   ;
13'd4192:weight<=16'b1111111110001110   ;
13'd4193:weight<=16'b0000000011010001   ;
13'd4194:weight<=16'b1111111111001010   ;
13'd4195:weight<=16'b1111111110011011   ;
13'd4196:weight<=16'b1111111110011110   ;
13'd4197:weight<=16'b0000000000000100   ;
13'd4198:weight<=16'b0000000010111010   ;
13'd4199:weight<=16'b0000000001010001   ;
13'd4200:weight<=16'b0000000111000101   ;
13'd4201:weight<=16'b0000000100111010   ;
13'd4202:weight<=16'b0000000001111110   ;
13'd4203:weight<=16'b0000000010100001   ;
13'd4204:weight<=16'b1111111111010000   ;
13'd4205:weight<=16'b1111111110110101   ;
13'd4206:weight<=16'b1111111010001101   ;
13'd4207:weight<=16'b1111111010010110   ;
13'd4208:weight<=16'b0000000010111110   ;
13'd4209:weight<=16'b1111111011111001   ;
13'd4210:weight<=16'b0000000000110101   ;
13'd4211:weight<=16'b1111111110010101   ;
13'd4212:weight<=16'b0000000000100110   ;
13'd4213:weight<=16'b1111111111010000   ;
13'd4214:weight<=16'b0000000001111011   ;
13'd4215:weight<=16'b1111111111110001   ;
13'd4216:weight<=16'b1111111100001011   ;
13'd4217:weight<=16'b0000000010000110   ;
13'd4218:weight<=16'b0000000010100010   ;
13'd4219:weight<=16'b1111111111101000   ;
13'd4220:weight<=16'b1111111111101110   ;
13'd4221:weight<=16'b1111111111011110   ;
13'd4222:weight<=16'b1111111111011100   ;
13'd4223:weight<=16'b0000000000000101   ;
13'd4224:weight<=16'b1111111111100001   ;
13'd4225:weight<=16'b1111111110100111   ;
13'd4226:weight<=16'b0000000001000110   ;
13'd4227:weight<=16'b0000000001101110   ;
13'd4228:weight<=16'b0000000000110010   ;
13'd4229:weight<=16'b0000000000110001   ;
13'd4230:weight<=16'b0000000000000011   ;
13'd4231:weight<=16'b0000000000001011   ;
13'd4232:weight<=16'b1111111110100100   ;
13'd4233:weight<=16'b1111111101011100   ;
13'd4234:weight<=16'b0000000000111100   ;
13'd4235:weight<=16'b0000000000010000   ;
13'd4236:weight<=16'b0000000001101000   ;
13'd4237:weight<=16'b0000000001000010   ;
13'd4238:weight<=16'b0000000010011001   ;
13'd4239:weight<=16'b1111111101100011   ;
13'd4240:weight<=16'b1111111110100101   ;
13'd4241:weight<=16'b1111111001100100   ;
13'd4242:weight<=16'b1111111111010100   ;
13'd4243:weight<=16'b1111111110110101   ;
13'd4244:weight<=16'b0000001001110000   ;
13'd4245:weight<=16'b0000000001000111   ;
13'd4246:weight<=16'b1111111101100110   ;
13'd4247:weight<=16'b0000000010111010   ;
13'd4248:weight<=16'b1111111111010110   ;
13'd4249:weight<=16'b0000000001010111   ;
13'd4250:weight<=16'b0000000111000101   ;
13'd4251:weight<=16'b0000000100111010   ;
13'd4252:weight<=16'b0000000001111110   ;
13'd4253:weight<=16'b0000000010100001   ;
13'd4254:weight<=16'b1111111111010000   ;
13'd4255:weight<=16'b1111111110110101   ;
13'd4256:weight<=16'b1111111010001101   ;
13'd4257:weight<=16'b1111111010010110   ;
13'd4258:weight<=16'b0000000010111110   ;
13'd4259:weight<=16'b1111111011111001   ;
13'd4260:weight<=16'b1111111111110011   ;
13'd4261:weight<=16'b1111111111000010   ;
13'd4262:weight<=16'b1111111111111110   ;
13'd4263:weight<=16'b0000000000011001   ;
13'd4264:weight<=16'b0000000000101000   ;
13'd4265:weight<=16'b1111111110110010   ;
13'd4266:weight<=16'b1111111111100111   ;
13'd4267:weight<=16'b0000000000000111   ;
13'd4268:weight<=16'b0000000000101010   ;
13'd4269:weight<=16'b0000000001000000   ;
13'd4270:weight<=16'b1111111111101110   ;
13'd4271:weight<=16'b1111111111011110   ;
13'd4272:weight<=16'b1111111111011100  ;
13'd4273:weight<=16'b0000000000000101   ;
13'd4274:weight<=16'b1111111111100001   ;
13'd4275:weight<=16'b1111111110100111   ;
13'd4276:weight<=16'b0000000001000110   ;
13'd4277:weight<=16'b0000000001101110   ;
13'd4278:weight<=16'b0000000000110010   ;
13'd4279:weight<=16'b0000000000110001   ;
13'd4280:weight<=16'b1111111101110110   ;
13'd4281:weight<=16'b0000000000100110   ;
13'd4282:weight<=16'b0000000100010001   ;
13'd4283:weight<=16'b0000000001000111   ;
13'd4284:weight<=16'b1111110111101101   ;
13'd4285:weight<=16'b0000000110010110   ;
13'd4286:weight<=16'b0000000000001000   ;
13'd4287:weight<=16'b0000000000100010   ;
13'd4288:weight<=16'b0000000001010111   ;
13'd4289:weight<=16'b1111111111101000   ;
13'd4290:weight<=16'b1111111110100101   ;
13'd4291:weight<=16'b1111111001100100   ;
13'd4292:weight<=16'b1111111111010100   ;
13'd4293:weight<=16'b1111111110110101   ;
13'd4294:weight<=16'b0000001001110000   ;
13'd4295:weight<=16'b0000000001000111   ;
13'd4296:weight<=16'b1111111101100110   ;
13'd4297:weight<=16'b0000000010111010   ;
13'd4298:weight<=16'b1111111111010110   ;
13'd4299:weight<=16'b0000000001010111   ;
13'd4300:weight<=16'b0000000001100110   ;
13'd4301:weight<=16'b0000000000110011   ;
13'd4302:weight<=16'b0000000001000110   ;
13'd4303:weight<=16'b1111111110001110   ;
13'd4304:weight<=16'b0000000000000101   ;
13'd4305:weight<=16'b1111111101110110   ;
13'd4306:weight<=16'b1111111110011110   ;
13'd4307:weight<=16'b1111111111011001   ;
13'd4308:weight<=16'b0000000001001110   ;
13'd4309:weight<=16'b0000000001101011   ;
13'd4310:weight<=16'b1111111111110011   ;
13'd4311:weight<=16'b1111111111000010   ;
13'd4312:weight<=16'b1111111111111110   ;
13'd4313:weight<=16'b0000000000011001   ;
13'd4314:weight<=16'b0000000000101000   ;
13'd4315:weight<=16'b1111111110110010   ;
13'd4316:weight<=16'b1111111111100111   ;
13'd4317:weight<=16'b0000000000000111   ;
13'd4318:weight<=16'b0000000000101010   ;
13'd4319:weight<=16'b0000000001000000   ;
13'd4320:weight<=16'b0000000000111101   ;
13'd4321:weight<=16'b1111111111001010   ;
13'd4322:weight<=16'b1111111110110110   ;
13'd4323:weight<=16'b0000000000010010   ;
13'd4324:weight<=16'b1111111111101000   ;
13'd4325:weight<=16'b1111111110001110   ;
13'd4326:weight<=16'b0000000000101000   ;
13'd4327:weight<=16'b0000000000100011   ;
13'd4328:weight<=16'b0000000001110100   ;
13'd4329:weight<=16'b0000000000000001   ;
13'd4330:weight<=16'b1111111101110110   ;
13'd4331:weight<=16'b0000000000100110   ;
13'd4332:weight<=16'b0000000100010001   ;
13'd4333:weight<=16'b0000000001000111   ;
13'd4334:weight<=16'b1111110111101101   ;
13'd4335:weight<=16'b0000000110010110   ;
13'd4336:weight<=16'b0000000000001000   ;
13'd4337:weight<=16'b0000000000100010   ;
13'd4338:weight<=16'b0000000001010111   ;
13'd4339:weight<=16'b1111111111101000   ;
13'd4340:weight<=16'b1111111101001101   ;
13'd4341:weight<=16'b1111111100011000   ;
13'd4342:weight<=16'b0000000110101010   ;
13'd4343:weight<=16'b1111111101111011   ;
13'd4344:weight<=16'b0000000001001000   ;
13'd4345:weight<=16'b0000000101110011   ;
13'd4346:weight<=16'b0000000100011101   ;
13'd4347:weight<=16'b1111111111100100   ;
13'd4348:weight<=16'b1111111011100110   ;
13'd4349:weight<=16'b1111111110010110   ;
13'd4350:weight<=16'b0000000001100110   ;
13'd4351:weight<=16'b0000000000110011   ;
13'd4352:weight<=16'b0000000001000110   ;
13'd4353:weight<=16'b1111111110001110   ;
13'd4354:weight<=16'b0000000000000101   ;
13'd4355:weight<=16'b1111111101110110   ;
13'd4356:weight<=16'b1111111110011110   ;
13'd4357:weight<=16'b1111111111011001   ;
13'd4358:weight<=16'b0000000001001110   ;
13'd4359:weight<=16'b0000000001101011   ;
13'd4360:weight<=16'b0000000001100000   ;
13'd4361:weight<=16'b0000000001101011   ;
13'd4362:weight<=16'b0000000000011101   ;
13'd4363:weight<=16'b1111111101101010   ;
13'd4364:weight<=16'b1111111101011100   ;
13'd4365:weight<=16'b0000000001101100   ;
13'd4366:weight<=16'b0000000000001000   ;
13'd4367:weight<=16'b0000000010001111   ;
13'd4368:weight<=16'b1111111110011011   ;
13'd4369:weight<=16'b1111111111110010   ;
13'd4370:weight<=16'b0000000000111101   ;
13'd4371:weight<=16'b1111111111001010   ;
13'd4372:weight<=16'b1111111110110110   ;
13'd4373:weight<=16'b0000000000010010   ;
13'd4374:weight<=16'b1111111111101000   ;
13'd4375:weight<=16'b1111111110001110   ;
13'd4376:weight<=16'b0000000000101000   ;
13'd4377:weight<=16'b0000000000100011   ;
13'd4378:weight<=16'b0000000001110100   ;
13'd4379:weight<=16'b0000000000000001   ;
13'd4380:weight<=16'b0000000000000101   ;
13'd4381:weight<=16'b0000000000101110   ;
13'd4382:weight<=16'b0000000000110001   ;
13'd4383:weight<=16'b1111111111100001   ;
13'd4384:weight<=16'b0000000001101110   ;
13'd4385:weight<=16'b1111111110111011   ;
13'd4386:weight<=16'b1111111111011010   ;
13'd4387:weight<=16'b1111111111000101   ;
13'd4388:weight<=16'b1111111110111011   ;
13'd4389:weight<=16'b0000000001010111   ;
13'd4390:weight<=16'b1111111101001101   ;
13'd4391:weight<=16'b1111111100011000   ;
13'd4392:weight<=16'b0000000110101010   ;
13'd4393:weight<=16'b1111111101111011   ;
13'd4394:weight<=16'b0000000001001000   ;
13'd4395:weight<=16'b0000000101110011   ;
13'd4396:weight<=16'b0000000100011101   ;
13'd4397:weight<=16'b1111111111100100   ;
13'd4398:weight<=16'b1111111011100110   ;
13'd4399:weight<=16'b1111111110010110   ;
13'd4400:weight<=16'b0000000000011010   ;
13'd4401:weight<=16'b1111111111010100   ;
13'd4402:weight<=16'b1111111111100001   ;
13'd4403:weight<=16'b1111111111101011   ;
13'd4404:weight<=16'b1111111111001010   ;
13'd4405:weight<=16'b1111111111011110   ;
13'd4406:weight<=16'b1111111111110000   ;
13'd4407:weight<=16'b0000000010011010   ;
13'd4408:weight<=16'b0000000001101011   ;
13'd4409:weight<=16'b1111111110111101   ;
13'd4410:weight<=16'b0000000001100000   ;
13'd4411:weight<=16'b0000000001101011   ;
13'd4412:weight<=16'b0000000000011101   ;
13'd4413:weight<=16'b1111111101101010   ;
13'd4414:weight<=16'b1111111101011100   ;
13'd4415:weight<=16'b0000000001101100   ;
13'd4416:weight<=16'b0000000000001000   ;
13'd4417:weight<=16'b0000000010001111   ;
13'd4418:weight<=16'b1111111110011011   ;
13'd4419:weight<=16'b1111111111110010   ;
13'd4420:weight<=16'b1111111111011010   ;
13'd4421:weight<=16'b0000000011110011   ;
13'd4422:weight<=16'b1111111101101011   ;
13'd4423:weight<=16'b1111111100000111   ;
13'd4424:weight<=16'b1111111110011011   ;
13'd4425:weight<=16'b1111111101111111   ;
13'd4426:weight<=16'b0000000001111010   ;
13'd4427:weight<=16'b0000000010001001   ;
13'd4428:weight<=16'b1111111110111000   ;
13'd4429:weight<=16'b0000000100110110   ;
13'd4430:weight<=16'b0000000000000101   ;
13'd4431:weight<=16'b0000000000101110   ;
13'd4432:weight<=16'b0000000000110001   ;
13'd4433:weight<=16'b1111111111100001   ;
13'd4434:weight<=16'b0000000001101110   ;
13'd4435:weight<=16'b1111111110111011   ;
13'd4436:weight<=16'b1111111111011010   ;
13'd4437:weight<=16'b1111111111000101   ;
13'd4438:weight<=16'b1111111110111011   ;
13'd4439:weight<=16'b0000000001010111   ;
13'd4440:weight<=16'b1111111111100011   ;
13'd4441:weight<=16'b0000000000000111   ;
13'd4442:weight<=16'b0000000001011110   ;
13'd4443:weight<=16'b0000000010011001   ;
13'd4444:weight<=16'b1111111111010001   ;
13'd4445:weight<=16'b0000000000011100   ;
13'd4446:weight<=16'b0000000000011001   ;
13'd4447:weight<=16'b0000000000100011   ;
13'd4448:weight<=16'b0000000001000111   ;
13'd4449:weight<=16'b1111111011101001   ;
13'd4450:weight<=16'b0000000000011010   ;
13'd4451:weight<=16'b1111111111010100   ;
13'd4452:weight<=16'b1111111111100001   ;
13'd4453:weight<=16'b1111111111101011   ;
13'd4454:weight<=16'b1111111111001010   ;
13'd4455:weight<=16'b1111111111011110   ;
13'd4456:weight<=16'b1111111111110000   ;
13'd4457:weight<=16'b0000000010011010   ;
13'd4458:weight<=16'b0000000001101011   ;
13'd4459:weight<=16'b1111111110111101   ;
13'd4460:weight<=16'b0000000000010000   ;
13'd4461:weight<=16'b1111111110000100   ;
13'd4462:weight<=16'b0000000001001011   ;
13'd4463:weight<=16'b1111111101111010   ;
13'd4464:weight<=16'b0000000000001101   ;
13'd4465:weight<=16'b0000000000010111   ;
13'd4466:weight<=16'b1111111111101101   ;
13'd4467:weight<=16'b0000000010001001   ;
13'd4468:weight<=16'b1111111111111100   ;
13'd4469:weight<=16'b0000000000100001   ;
13'd4470:weight<=16'b1111111111011010   ;
13'd4471:weight<=16'b0000000011110011   ;
13'd4472:weight<=16'b1111111101101011   ;
13'd4473:weight<=16'b1111111100000111   ;
13'd4474:weight<=16'b1111111110011011   ;
13'd4475:weight<=16'b1111111101111111   ;
13'd4476:weight<=16'b0000000001111010   ;
13'd4477:weight<=16'b0000000010001001   ;
13'd4478:weight<=16'b1111111110111000   ;
13'd4479:weight<=16'b0000000100110110   ;
13'd4480:weight<=16'b0000000001011001   ;
13'd4481:weight<=16'b1111111111010101   ;
13'd4482:weight<=16'b1111111111101100   ;
13'd4483:weight<=16'b1111111111111110   ;
13'd4484:weight<=16'b0000000100101101   ;
13'd4485:weight<=16'b1111111111001001   ;
13'd4486:weight<=16'b1111111101011010   ;
13'd4487:weight<=16'b1111111101111111   ;
13'd4488:weight<=16'b1111111100111110   ;
13'd4489:weight<=16'b0000000100100000   ;
13'd4490:weight<=16'b1111111111100011   ;
13'd4491:weight<=16'b0000000000000111   ;
13'd4492:weight<=16'b0000000001011110   ;
13'd4493:weight<=16'b0000000010011001   ;
13'd4494:weight<=16'b1111111111010001   ;
13'd4495:weight<=16'b0000000000011100   ;
13'd4496:weight<=16'b0000000000011001   ;
13'd4497:weight<=16'b0000000000100011   ;
13'd4498:weight<=16'b0000000001000111   ;
13'd4499:weight<=16'b1111111011101001   ;
13'd4500:weight<=16'b0000000001011101   ;
13'd4501:weight<=16'b1111111111111110   ;
13'd4502:weight<=16'b1111111111000011   ;
13'd4503:weight<=16'b0000000001010110   ;
13'd4504:weight<=16'b1111111110100011   ;
13'd4505:weight<=16'b0000000000110001   ;
13'd4506:weight<=16'b0000000000001001   ;
13'd4507:weight<=16'b0000000000001101   ;
13'd4508:weight<=16'b1111111111000010   ;
13'd4509:weight<=16'b1111111111010000   ;
13'd4510:weight<=16'b0000000000010000   ;
13'd4511:weight<=16'b1111111110000100   ;
13'd4512:weight<=16'b0000000001001011   ;
13'd4513:weight<=16'b1111111101111010   ;
13'd4514:weight<=16'b0000000000001101   ;
13'd4515:weight<=16'b0000000000010111   ;
13'd4516:weight<=16'b1111111111101101   ;
13'd4517:weight<=16'b0000000010001001   ;
13'd4518:weight<=16'b1111111111111100   ;
13'd4519:weight<=16'b0000000000100001   ;
13'd4520:weight<=16'b0000000001011110   ;
13'd4521:weight<=16'b0000000111101110   ;
13'd4522:weight<=16'b1111111111111001   ;
13'd4523:weight<=16'b0000000000001100   ;
13'd4524:weight<=16'b1111111101100110   ;
13'd4525:weight<=16'b1111111101111101   ;
13'd4526:weight<=16'b1111111110001101   ;
13'd4527:weight<=16'b1111111100101010   ;
13'd4528:weight<=16'b0000000001110110   ;
13'd4529:weight<=16'b1111111111011000   ;
13'd4530:weight<=16'b0000000001011001   ;
13'd4531:weight<=16'b1111111111010101   ;
13'd4532:weight<=16'b1111111111101100   ;
13'd4533:weight<=16'b1111111111111110   ;
13'd4534:weight<=16'b0000000100101101   ;
13'd4535:weight<=16'b1111111111001001   ;
13'd4536:weight<=16'b1111111101011010   ;
13'd4537:weight<=16'b1111111101111111   ;
13'd4538:weight<=16'b1111111100111110   ;
13'd4539:weight<=16'b0000000100100000   ;
13'd4540:weight<=16'b0000000001101111   ;
13'd4541:weight<=16'b1111111111111011   ;
13'd4542:weight<=16'b0000000001111110   ;
13'd4543:weight<=16'b1111111100111110   ;
13'd4544:weight<=16'b0000000001101001   ;
13'd4545:weight<=16'b1111111111110001   ;
13'd4546:weight<=16'b1111111110101110   ;
13'd4547:weight<=16'b0000000011000010   ;
13'd4548:weight<=16'b1111111101010110   ;
13'd4549:weight<=16'b0000000000000110   ;
13'd4550:weight<=16'b0000000001011101   ;
13'd4551:weight<=16'b1111111111111110   ;
13'd4552:weight<=16'b1111111111000011   ;
13'd4553:weight<=16'b0000000001010110   ;
13'd4554:weight<=16'b1111111110100011   ;
13'd4555:weight<=16'b0000000000110001   ;
13'd4556:weight<=16'b0000000000001001   ;
13'd4557:weight<=16'b0000000000001101   ;
13'd4558:weight<=16'b1111111111000010   ;
13'd4559:weight<=16'b1111111111010000   ;
13'd4560:weight<=16'b0000000000110101   ;
13'd4561:weight<=16'b0000000010011011   ;
13'd4562:weight<=16'b0000000000000001   ;
13'd4563:weight<=16'b1111111110011101   ;
13'd4564:weight<=16'b0000000000011000   ;
13'd4565:weight<=16'b0000000110011100   ;
13'd4566:weight<=16'b1111111100100101   ;
13'd4567:weight<=16'b1111111111010010   ;
13'd4568:weight<=16'b1111111111011010   ;
13'd4569:weight<=16'b1111111101011000   ;
13'd4570:weight<=16'b0000000001011110   ;
13'd4571:weight<=16'b0000000111101110   ;
13'd4572:weight<=16'b1111111111111001   ;
13'd4573:weight<=16'b0000000000001100   ;
13'd4574:weight<=16'b1111111101100110   ;
13'd4575:weight<=16'b1111111101111101   ;
13'd4576:weight<=16'b1111111110001101   ;
13'd4577:weight<=16'b1111111100101010   ;
13'd4578:weight<=16'b0000000001110110   ;
13'd4579:weight<=16'b1111111111011000   ;
13'd4580:weight<=16'b1111111111101010   ;
13'd4581:weight<=16'b1111111111110111   ;
13'd4582:weight<=16'b0000000010001111   ;
13'd4583:weight<=16'b0000000000000011   ;
13'd4584:weight<=16'b0000000010001110   ;
13'd4585:weight<=16'b0000000001001010   ;
13'd4586:weight<=16'b1111111111000111   ;
13'd4587:weight<=16'b1111111111100010   ;
13'd4588:weight<=16'b1111111101001110   ;
13'd4589:weight<=16'b0000000000000010   ;
13'd4590:weight<=16'b0000000001101111   ;
13'd4591:weight<=16'b1111111111111011   ;
13'd4592:weight<=16'b0000000001111110   ;
13'd4593:weight<=16'b1111111100111110   ;
13'd4594:weight<=16'b0000000001101001   ;
13'd4595:weight<=16'b1111111111110001   ;
13'd4596:weight<=16'b1111111110101110   ;
13'd4597:weight<=16'b0000000011000010   ;
13'd4598:weight<=16'b1111111101010110   ;
13'd4599:weight<=16'b0000000000000110   ;
13'd4600:weight<=16'b0000000000011011   ;
13'd4601:weight<=16'b0000000011000010   ;
13'd4602:weight<=16'b1111111101101100   ;
13'd4603:weight<=16'b0000000001100000   ;
13'd4604:weight<=16'b0000000001000100   ;
13'd4605:weight<=16'b1111111110101111   ;
13'd4606:weight<=16'b1111111111100000   ;
13'd4607:weight<=16'b1111111111100100   ;
13'd4608:weight<=16'b0000000000101000   ;
13'd4609:weight<=16'b1111111110010101   ;
13'd4610:weight<=16'b0000000000110101   ;
13'd4611:weight<=16'b0000000010011011   ;
13'd4612:weight<=16'b0000000000000001   ;
13'd4613:weight<=16'b1111111110011101   ;
13'd4614:weight<=16'b0000000000011000   ;
13'd4615:weight<=16'b0000000110011100   ;
13'd4616:weight<=16'b1111111100100101   ;
13'd4617:weight<=16'b1111111111010010   ;
13'd4618:weight<=16'b1111111111011010   ;
13'd4619:weight<=16'b1111111101011000   ;
13'd4620:weight<=16'b0000000011010010   ;
13'd4621:weight<=16'b0000000000100011   ;
13'd4622:weight<=16'b0000000000010010   ;
13'd4623:weight<=16'b1111111010111011   ;
13'd4624:weight<=16'b0000000000000100   ;
13'd4625:weight<=16'b0000000011010111   ;
13'd4626:weight<=16'b1111111011110000   ;
13'd4627:weight<=16'b0000000001001101   ;
13'd4628:weight<=16'b0000000011010010   ;
13'd4629:weight<=16'b1111111101111000   ;
13'd4630:weight<=16'b1111111111101010   ;
13'd4631:weight<=16'b1111111111110111   ;
13'd4632:weight<=16'b0000000010001111   ;
13'd4633:weight<=16'b0000000000000011   ;
13'd4634:weight<=16'b0000000010001110   ;
13'd4635:weight<=16'b0000000001001010   ;
13'd4636:weight<=16'b1111111111000111   ;
13'd4637:weight<=16'b1111111111100010   ;
13'd4638:weight<=16'b1111111101001110   ;
13'd4639:weight<=16'b0000000000000010   ;
13'd4640:weight<=16'b0000000000100111   ;
13'd4641:weight<=16'b0000000001011000   ;
13'd4642:weight<=16'b0000000000001101   ;
13'd4643:weight<=16'b1111111110000111   ;
13'd4644:weight<=16'b0000000001110000   ;
13'd4645:weight<=16'b0000000000011000   ;
13'd4646:weight<=16'b1111111111010011   ;
13'd4647:weight<=16'b1111111101100001   ;
13'd4648:weight<=16'b0000000100000010   ;
13'd4649:weight<=16'b1111111101100011   ;
13'd4650:weight<=16'b0000000000011011   ;
13'd4651:weight<=16'b0000000011000010   ;
13'd4652:weight<=16'b1111111101101100   ;
13'd4653:weight<=16'b0000000001100000   ;
13'd4654:weight<=16'b0000000001000100   ;
13'd4655:weight<=16'b1111111110101111   ;
13'd4656:weight<=16'b1111111111100000   ;
13'd4657:weight<=16'b1111111111100100   ;
13'd4658:weight<=16'b0000000000101000   ;
13'd4659:weight<=16'b1111111110010101   ;
13'd4660:weight<=16'b0000000010000110   ;
13'd4661:weight<=16'b0000000001111111   ;
13'd4662:weight<=16'b1111111111100000   ;
13'd4663:weight<=16'b1111111100111101   ;
13'd4664:weight<=16'b1111111111111010   ;
13'd4665:weight<=16'b1111111111001101   ;
13'd4666:weight<=16'b1111111110001011   ;
13'd4667:weight<=16'b0000000010011100   ;
13'd4668:weight<=16'b0000000011010011   ;
13'd4669:weight<=16'b1111111100100100   ;
13'd4670:weight<=16'b0000000011010010   ;
13'd4671:weight<=16'b0000000000100011   ;
13'd4672:weight<=16'b0000000000010010   ;
13'd4673:weight<=16'b1111111010111011   ;
13'd4674:weight<=16'b0000000000000100   ;
13'd4675:weight<=16'b0000000011010111   ;
13'd4676:weight<=16'b1111111011110000   ;
13'd4677:weight<=16'b0000000001001101   ;
13'd4678:weight<=16'b0000000011010010   ;
13'd4679:weight<=16'b1111111101111000   ;
13'd4680:weight<=16'b0000000000000101   ;
13'd4681:weight<=16'b0000000011111011   ;
13'd4682:weight<=16'b1111111111101010   ;
13'd4683:weight<=16'b1111111110010010   ;
13'd4684:weight<=16'b1111111111111001   ;
13'd4685:weight<=16'b0000000001011111   ;
13'd4686:weight<=16'b0000000000001000   ;
13'd4687:weight<=16'b1111111101100111   ;
13'd4688:weight<=16'b0000000001110000   ;
13'd4689:weight<=16'b1111111101111010   ;
13'd4690:weight<=16'b0000000000100111   ;
13'd4691:weight<=16'b0000000001011000   ;
13'd4692:weight<=16'b0000000000001101   ;
13'd4693:weight<=16'b1111111110000111   ;
13'd4694:weight<=16'b0000000001110000   ;
13'd4695:weight<=16'b0000000000011000   ;
13'd4696:weight<=16'b1111111111010011   ;
13'd4697:weight<=16'b1111111101100001   ;
13'd4698:weight<=16'b0000000100000010   ;
13'd4699:weight<=16'b1111111101100011   ;
13'd4700:weight<=16'b1111111110011001   ;
13'd4701:weight<=16'b1111111111011100   ;
13'd4702:weight<=16'b1111111110011000   ;
13'd4703:weight<=16'b0000000001010111   ;
13'd4704:weight<=16'b0000000010111001   ;
13'd4705:weight<=16'b0000000001000101   ;
13'd4706:weight<=16'b0000000000001010   ;
13'd4707:weight<=16'b1111111110010110   ;
13'd4708:weight<=16'b0000000001111111   ;
13'd4709:weight<=16'b1111111111001011   ;
13'd4710:weight<=16'b0000000010000110   ;
13'd4711:weight<=16'b0000000001111111   ;
13'd4712:weight<=16'b1111111111100000   ;
13'd4713:weight<=16'b1111111100111101   ;
13'd4714:weight<=16'b1111111111111010   ;
13'd4715:weight<=16'b1111111111001101   ;
13'd4716:weight<=16'b1111111110001011   ;
13'd4717:weight<=16'b0000000010011100   ;
13'd4718:weight<=16'b0000000011010011   ;
13'd4719:weight<=16'b1111111100100100  ;
13'd4720:weight<=16'b1111111101000101   ;
13'd4721:weight<=16'b0000000010010010   ;
13'd4722:weight<=16'b0000000011001011   ;
13'd4723:weight<=16'b0000000001011111   ;
13'd4724:weight<=16'b0000000100001011   ;
13'd4725:weight<=16'b1111111111000100   ;
13'd4726:weight<=16'b1111111111000010   ;
13'd4727:weight<=16'b1111111100110011   ;
13'd4728:weight<=16'b1111111111100111   ;
13'd4729:weight<=16'b1111111110100100   ;
13'd4730:weight<=16'b0000000000000101   ;
13'd4731:weight<=16'b0000000011111011   ;
13'd4732:weight<=16'b1111111111101010   ;
13'd4733:weight<=16'b1111111110010010   ;
13'd4734:weight<=16'b1111111111111001   ;
13'd4735:weight<=16'b0000000001011111   ;
13'd4736:weight<=16'b0000000000001000   ;
13'd4737:weight<=16'b1111111101100111   ;
13'd4738:weight<=16'b0000000001110000   ;
13'd4739:weight<=16'b1111111101111010   ;
13'd4740:weight<=16'b0000000001010111   ;
13'd4741:weight<=16'b0000000001111011   ;
13'd4742:weight<=16'b0000000000110111   ;
13'd4743:weight<=16'b0000000000110000   ;
13'd4744:weight<=16'b1111111111000010   ;
13'd4745:weight<=16'b1111111111000000   ;
13'd4746:weight<=16'b0000000001101010   ;
13'd4747:weight<=16'b1111111110110110   ;
13'd4748:weight<=16'b1111111100000010   ;
13'd4749:weight<=16'b0000000001000110   ;
13'd4750:weight<=16'b1111111110011001   ;
13'd4751:weight<=16'b1111111111011100   ;
13'd4752:weight<=16'b1111111110011000   ;
13'd4753:weight<=16'b0000000001010111   ;
13'd4754:weight<=16'b0000000010111001   ;
13'd4755:weight<=16'b0000000001000101   ;
13'd4756:weight<=16'b0000000000001010   ;
13'd4757:weight<=16'b1111111110010110   ;
13'd4758:weight<=16'b0000000001111111   ;
13'd4759:weight<=16'b1111111111001011   ;
13'd4760:weight<=16'b1111111111001000   ;
13'd4761:weight<=16'b1111111111101110   ;
13'd4762:weight<=16'b0000000010001110   ;
13'd4763:weight<=16'b1111111111110111   ;
13'd4764:weight<=16'b0000000000011110   ;
13'd4765:weight<=16'b1111111111101110   ;
13'd4766:weight<=16'b0000000001000011   ;
13'd4767:weight<=16'b0000000000011101   ;
13'd4768:weight<=16'b1111111111010101   ;
13'd4769:weight<=16'b1111111111001011   ;
13'd4770:weight<=16'b1111111101000101   ;
13'd4771:weight<=16'b0000000010010010   ;
13'd4772:weight<=16'b0000000011001011   ;
13'd4773:weight<=16'b0000000001011111   ;
13'd4774:weight<=16'b0000000100001011   ;
13'd4775:weight<=16'b1111111111000100   ;
13'd4776:weight<=16'b1111111111000010   ;
13'd4777:weight<=16'b1111111100110011   ;
13'd4778:weight<=16'b1111111111100111   ;
13'd4779:weight<=16'b1111111110100100   ;
13'd4780:weight<=16'b1111111110101100   ;
13'd4781:weight<=16'b1111111110100111   ;
13'd4782:weight<=16'b0000000001100100   ;
13'd4783:weight<=16'b0000000000010001   ;
13'd4784:weight<=16'b1111111111101001   ;
13'd4785:weight<=16'b1111111111010100   ;
13'd4786:weight<=16'b0000000000111010   ;
13'd4787:weight<=16'b1111111111101111   ;
13'd4788:weight<=16'b0000000001000000   ;
13'd4789:weight<=16'b0000000000000001   ;
13'd4790:weight<=16'b0000000001010111   ;
13'd4791:weight<=16'b0000000001111011   ;
13'd4792:weight<=16'b0000000000110111   ;
13'd4793:weight<=16'b0000000000110000   ;
13'd4794:weight<=16'b1111111111000010   ;
13'd4795:weight<=16'b1111111111000000   ;
13'd4796:weight<=16'b0000000001101010   ;
13'd4797:weight<=16'b1111111110110110   ;
13'd4798:weight<=16'b1111111100000010   ;
13'd4799:weight<=16'b0000000001000110   ;
13'd4800:weight<=16'b1111111111101100   ;
13'd4801:weight<=16'b0000000001011101   ;
13'd4802:weight<=16'b1111111111110010   ;
13'd4803:weight<=16'b1111111111011101   ;
13'd4804:weight<=16'b0000000001000010   ;
13'd4805:weight<=16'b1111111111110111   ;
13'd4806:weight<=16'b0000000000000011   ;
13'd4807:weight<=16'b0000000000000000   ;
13'd4808:weight<=16'b1111111111001100   ;
13'd4809:weight<=16'b0000000000001100   ;
13'd4810:weight<=16'b1111111111001000   ;
13'd4811:weight<=16'b1111111111101110   ;
13'd4812:weight<=16'b0000000010001110   ;
13'd4813:weight<=16'b1111111111110111   ;
13'd4814:weight<=16'b0000000000011110   ;
13'd4815:weight<=16'b1111111111101110   ;
13'd4816:weight<=16'b0000000001000011   ;
13'd4817:weight<=16'b0000000000011101   ;
13'd4818:weight<=16'b1111111111010101   ;
13'd4819:weight<=16'b1111111111001011   ;
13'd4820:weight<=16'b1111111111111000   ;
13'd4821:weight<=16'b0000000101011111   ;
13'd4822:weight<=16'b1111111101110011   ;
13'd4823:weight<=16'b1111111110010010   ;
13'd4824:weight<=16'b1111111101110101   ;
13'd4825:weight<=16'b1111111111001000   ;
13'd4826:weight<=16'b0000000001010111   ;
13'd4827:weight<=16'b0000000011100000   ;
13'd4828:weight<=16'b0000000000011100   ;
13'd4829:weight<=16'b1111111100110111   ;
13'd4830:weight<=16'b1111111110101100   ;
13'd4831:weight<=16'b1111111110100111   ;
13'd4832:weight<=16'b0000000001100100   ;
13'd4833:weight<=16'b0000000000010001   ;
13'd4834:weight<=16'b1111111111101001   ;
13'd4835:weight<=16'b1111111111010100   ;
13'd4836:weight<=16'b0000000000111010   ;
13'd4837:weight<=16'b1111111111101111   ;
13'd4838:weight<=16'b0000000001000000   ;
13'd4839:weight<=16'b0000000000000001   ;
13'd4840:weight<=16'b0000000000001010   ;
13'd4841:weight<=16'b1111111111110111   ;
13'd4842:weight<=16'b0000000000110010   ;
13'd4843:weight<=16'b0000000001001010   ;
13'd4844:weight<=16'b0000000000001011   ;
13'd4845:weight<=16'b0000000000110101   ;
13'd4846:weight<=16'b1111111111110011   ;
13'd4847:weight<=16'b0000000000110110   ;
13'd4848:weight<=16'b1111111110011001   ;
13'd4849:weight<=16'b1111111110110001   ;
13'd4850:weight<=16'b1111111111101100   ;
13'd4851:weight<=16'b0000000001011101   ;
13'd4852:weight<=16'b1111111111110010   ;
13'd4853:weight<=16'b1111111111011101   ;
13'd4854:weight<=16'b0000000001000010   ;
13'd4855:weight<=16'b1111111111110111   ;
13'd4856:weight<=16'b0000000000000011   ;
13'd4857:weight<=16'b0000000000000000   ;
13'd4858:weight<=16'b1111111111001100   ;
13'd4859:weight<=16'b0000000000001100   ;
13'd4860:weight<=16'b1111111111011110   ;
13'd4861:weight<=16'b1111111110011010   ;
13'd4862:weight<=16'b1111111110101010   ;
13'd4863:weight<=16'b0000000000100111   ;
13'd4864:weight<=16'b0000000010110000   ;
13'd4865:weight<=16'b0000000000101100   ;
13'd4866:weight<=16'b1111111111110101   ;
13'd4867:weight<=16'b0000000010000000   ;
13'd4868:weight<=16'b1111111111101101   ;
13'd4869:weight<=16'b1111111110001011   ;
13'd4870:weight<=16'b1111111111111000   ;
13'd4871:weight<=16'b0000000101011111   ;
13'd4872:weight<=16'b1111111101110011   ;
13'd4873:weight<=16'b1111111110010010   ;
13'd4874:weight<=16'b1111111101110101   ;
13'd4875:weight<=16'b1111111111001000   ;
13'd4876:weight<=16'b0000000001010111   ;
13'd4877:weight<=16'b0000000011100000   ;
13'd4878:weight<=16'b0000000000011100   ;
13'd4879:weight<=16'b1111111100110111   ;
13'd4880:weight<=16'b1111111110010011   ;
13'd4881:weight<=16'b1111111111001110   ;
13'd4882:weight<=16'b0000000010111110   ;
13'd4883:weight<=16'b1111111111001001   ;
13'd4884:weight<=16'b1111111111100000   ;
13'd4885:weight<=16'b0000000000000101   ;
13'd4886:weight<=16'b1111111110110111   ;
13'd4887:weight<=16'b0000000001101011   ;
13'd4888:weight<=16'b0000000000000100   ;
13'd4889:weight<=16'b0000000000110101   ;
13'd4890:weight<=16'b0000000000001010   ;
13'd4891:weight<=16'b1111111111110111   ;
13'd4892:weight<=16'b0000000000110010   ;
13'd4893:weight<=16'b0000000001001010   ;
13'd4894:weight<=16'b0000000000001011   ;
13'd4895:weight<=16'b0000000000110101   ;
13'd4896:weight<=16'b1111111111110011   ;
13'd4897:weight<=16'b0000000000110110   ;
13'd4898:weight<=16'b1111111110011001   ;
13'd4899:weight<=16'b1111111110110001   ;
13'd4900:weight<=16'b1111111110100010   ;
13'd4901:weight<=16'b1111111110101000   ;
13'd4902:weight<=16'b1111111111000001   ;
13'd4903:weight<=16'b0000000010100111   ;
13'd4904:weight<=16'b0000000000010100  ;
13'd4905:weight<=16'b0000000000010011   ;
13'd4906:weight<=16'b1111111110110100   ;
13'd4907:weight<=16'b0000000001101111   ;
13'd4908:weight<=16'b0000000001011011   ;
13'd4909:weight<=16'b1111111111100100   ;
13'd4910:weight<=16'b1111111111011110   ;
13'd4911:weight<=16'b1111111110011010   ;
13'd4912:weight<=16'b1111111110101010   ;
13'd4913:weight<=16'b0000000000100111   ;
13'd4914:weight<=16'b0000000010110000   ;
13'd4915:weight<=16'b0000000000101100   ;
13'd4916:weight<=16'b1111111111110101   ;
13'd4917:weight<=16'b0000000010000000   ;
13'd4918:weight<=16'b1111111111101101   ;
13'd4919:weight<=16'b1111111110001011   ;
13'd4920:weight<=16'b0000000010100111   ;
13'd4921:weight<=16'b1111111010111110   ;
13'd4922:weight<=16'b1111111110011110   ;
13'd4923:weight<=16'b0000000000001111   ;
13'd4924:weight<=16'b0000000000001111   ;
13'd4925:weight<=16'b0000000011101110   ;
13'd4926:weight<=16'b1111111111000000   ;
13'd4927:weight<=16'b1111111111001111   ;
13'd4928:weight<=16'b0000000010000100   ;
13'd4929:weight<=16'b0000000001111010   ;
13'd4930:weight<=16'b1111111110010011   ;
13'd4931:weight<=16'b1111111111001110   ;
13'd4932:weight<=16'b0000000010111110   ;
13'd4933:weight<=16'b1111111111001001   ;
13'd4934:weight<=16'b1111111111100000   ;
13'd4935:weight<=16'b0000000000000101   ;
13'd4936:weight<=16'b1111111110110111   ;
13'd4937:weight<=16'b0000000001101011   ;
13'd4938:weight<=16'b0000000000000100   ;
13'd4939:weight<=16'b0000000000110101   ;
13'd4940:weight<=16'b1111111110011110   ;
13'd4941:weight<=16'b0000000010010000   ;
13'd4942:weight<=16'b1111111111110111   ;
13'd4943:weight<=16'b0000000000100001   ;
13'd4944:weight<=16'b1111111110010101   ;
13'd4945:weight<=16'b0000000001011111   ;
13'd4946:weight<=16'b0000000000100100   ;
13'd4947:weight<=16'b1111111110111101   ;
13'd4948:weight<=16'b0000000000111110   ;
13'd4949:weight<=16'b1111111110111101   ;
13'd4950:weight<=16'b1111111110100010   ;
13'd4951:weight<=16'b1111111110101000   ;
13'd4952:weight<=16'b1111111111000001   ;
13'd4953:weight<=16'b0000000010100111   ;
13'd4954:weight<=16'b0000000000010100   ;
13'd4955:weight<=16'b0000000000010011   ;
13'd4956:weight<=16'b1111111110110100   ;
13'd4957:weight<=16'b0000000001101111   ;
13'd4958:weight<=16'b0000000001011011   ;
13'd4959:weight<=16'b1111111111100100   ;
13'd4960:weight<=16'b1111111110110011   ;
13'd4961:weight<=16'b0000000000000001   ;
13'd4962:weight<=16'b0000000000001001   ;
13'd4963:weight<=16'b0000000001000001   ;
13'd4964:weight<=16'b0000000000011010   ;
13'd4965:weight<=16'b0000000001101001   ;
13'd4966:weight<=16'b0000000000110101   ;
13'd4967:weight<=16'b1111111111001111   ;
13'd4968:weight<=16'b1111111110001110   ;
13'd4969:weight<=16'b1111111111100011   ;
13'd4970:weight<=16'b0000000010100111   ;
13'd4971:weight<=16'b1111111010111110   ;
13'd4972:weight<=16'b1111111110011110   ;
13'd4973:weight<=16'b0000000000001111   ;
13'd4974:weight<=16'b0000000000001111   ;
13'd4975:weight<=16'b0000000011101110   ;
13'd4976:weight<=16'b1111111111000000   ;
13'd4977:weight<=16'b1111111111001111   ;
13'd4978:weight<=16'b0000000010000100   ;
13'd4979:weight<=16'b0000000001111010   ;
13'd4980:weight<=16'b1111111111110111   ;
13'd4981:weight<=16'b0000000001011111   ;
13'd4982:weight<=16'b1111111110111011   ;
13'd4983:weight<=16'b0000000001110011   ;
13'd4984:weight<=16'b0000000000100000   ;
13'd4985:weight<=16'b0000000010010000   ;
13'd4986:weight<=16'b1111111111110101   ;
13'd4987:weight<=16'b0000000001100000   ;
13'd4988:weight<=16'b1111111101001000   ;
13'd4989:weight<=16'b1111111111001001   ;
13'd4990:weight<=16'b1111111110011110   ;
13'd4991:weight<=16'b0000000010010000   ;
13'd4992:weight<=16'b1111111111110111   ;
13'd4993:weight<=16'b0000000000100001   ;
13'd4994:weight<=16'b1111111110010101   ;
13'd4995:weight<=16'b0000000001011111   ;
13'd4996:weight<=16'b0000000000100100   ;
13'd4997:weight<=16'b1111111110111101   ;
13'd4998:weight<=16'b0000000000111110   ;
13'd4999:weight<=16'b1111111110111101   ;
13'd5000:weight<=16'b0000000001110101   ;
13'd5001:weight<=16'b1111111101111000   ;
13'd5002:weight<=16'b0000000000101110   ;
13'd5003:weight<=16'b0000000001111100   ;
13'd5004:weight<=16'b0000000001010100   ;
13'd5005:weight<=16'b0000000000001011   ;
13'd5006:weight<=16'b1111111111010111   ;
13'd5007:weight<=16'b0000000000111010   ;
13'd5008:weight<=16'b1111111110010101   ;
13'd5009:weight<=16'b1111111110010111   ;
13'd5010:weight<=16'b1111111110110011   ;
13'd5011:weight<=16'b0000000000000001   ;
13'd5012:weight<=16'b0000000000001001   ;
13'd5013:weight<=16'b0000000001000001   ;
13'd5014:weight<=16'b0000000000011010   ;
13'd5015:weight<=16'b0000000001101001   ;
13'd5016:weight<=16'b0000000000110101   ;
13'd5017:weight<=16'b1111111111001111   ;
13'd5018:weight<=16'b1111111110001110   ;
13'd5019:weight<=16'b1111111111100011   ;
13'd5020:weight<=16'b1111111111011000   ;
13'd5021:weight<=16'b0000000000100000   ;
13'd5022:weight<=16'b0000000000011100   ;
13'd5023:weight<=16'b1111111101111011   ;
13'd5024:weight<=16'b0000000010010010   ;
13'd5025:weight<=16'b0000000011010101   ;
13'd5026:weight<=16'b0000000000011001   ;
13'd5027:weight<=16'b1111111110001001   ;
13'd5028:weight<=16'b1111111110100110   ;
13'd5029:weight<=16'b1111111111100100   ;
13'd5030:weight<=16'b1111111111110111   ;
13'd5031:weight<=16'b0000000001011111   ;
13'd5032:weight<=16'b1111111110111011   ;
13'd5033:weight<=16'b0000000001110011   ;
13'd5034:weight<=16'b0000000000100000   ;
13'd5035:weight<=16'b0000000010010000   ;
13'd5036:weight<=16'b1111111111110101   ;
13'd5037:weight<=16'b0000000001100000   ;
13'd5038:weight<=16'b1111111101001000   ;
13'd5039:weight<=16'b1111111111001001   ;
13'd5040:weight<=16'b0000000000010101   ;
13'd5041:weight<=16'b1111111111000000   ;
13'd5042:weight<=16'b0000000011000010   ;
13'd5043:weight<=16'b0000000001100100   ;
13'd5044:weight<=16'b0000000010100011   ;
13'd5045:weight<=16'b0000000010100000   ;
13'd5046:weight<=16'b1111111110101011   ;
13'd5047:weight<=16'b1111111100101000   ;
13'd5048:weight<=16'b1111111110100010   ;
13'd5049:weight<=16'b1111111110100101   ;
13'd5050:weight<=16'b0000000001110101   ;
13'd5051:weight<=16'b1111111101111000   ;
13'd5052:weight<=16'b0000000000101110   ;
13'd5053:weight<=16'b0000000001111100   ;
13'd5054:weight<=16'b0000000001010100   ;
13'd5055:weight<=16'b0000000000001011   ;
13'd5056:weight<=16'b1111111111010111   ;
13'd5057:weight<=16'b0000000000111010   ;
13'd5058:weight<=16'b1111111110010101   ;
13'd5059:weight<=16'b1111111110010111   ;
13'd5060:weight<=16'b1111111110100000   ;
13'd5061:weight<=16'b1111111110111100   ;
13'd5062:weight<=16'b0000000010000001   ;
13'd5063:weight<=16'b0000000000001100   ;
13'd5064:weight<=16'b1111111110110100   ;
13'd5065:weight<=16'b0000000001100001   ;
13'd5066:weight<=16'b0000000010011101   ;
13'd5067:weight<=16'b1111111111110100   ;
13'd5068:weight<=16'b1111111110010011   ;
13'd5069:weight<=16'b0000000000001111   ;
13'd5070:weight<=16'b1111111111011000   ;
13'd5071:weight<=16'b0000000000100000   ;
13'd5072:weight<=16'b0000000000011100   ;
13'd5073:weight<=16'b1111111101111011   ;
13'd5074:weight<=16'b0000000010010010   ;
13'd5075:weight<=16'b0000000011010101   ;
13'd5076:weight<=16'b0000000000011001   ;
13'd5077:weight<=16'b1111111110001001   ;
13'd5078:weight<=16'b1111111110100110   ;
13'd5079:weight<=16'b1111111111100100   ;
13'd5080:weight<=16'b0000000000100101   ;
13'd5081:weight<=16'b0000000001111010   ;
13'd5082:weight<=16'b0000000010110111   ;
13'd5083:weight<=16'b1111111111000011   ;
13'd5084:weight<=16'b0000000000011010   ;
13'd5085:weight<=16'b1111111101110000   ;
13'd5086:weight<=16'b0000000101001101   ;
13'd5087:weight<=16'b1111111011011000   ;
13'd5088:weight<=16'b0000000001110001   ;
13'd5089:weight<=16'b1111111011010001   ;
13'd5090:weight<=16'b0000000000010101   ;
13'd5091:weight<=16'b1111111111000000   ;
13'd5092:weight<=16'b0000000011000010   ;
13'd5093:weight<=16'b0000000001100100   ;
13'd5094:weight<=16'b0000000010100011   ;
13'd5095:weight<=16'b0000000010100000   ;
13'd5096:weight<=16'b1111111110101011   ;
13'd5097:weight<=16'b1111111100101000   ;
13'd5098:weight<=16'b1111111110100010   ;
13'd5099:weight<=16'b1111111110100101   ;
13'd5100:weight<=16'b1111111100110010   ;
13'd5101:weight<=16'b0000001001111001   ;
13'd5102:weight<=16'b0000000110001110   ;
13'd5103:weight<=16'b1111111111110110   ;
13'd5104:weight<=16'b1111110111011011   ;
13'd5105:weight<=16'b0000000010000000   ;
13'd5106:weight<=16'b0000000000101000   ;
13'd5107:weight<=16'b1111111111000111   ;
13'd5108:weight<=16'b1111111010011111   ;
13'd5109:weight<=16'b0000000010000100   ;
13'd5110:weight<=16'b1111111110100000   ;
13'd5111:weight<=16'b1111111110111100   ;
13'd5112:weight<=16'b0000000010000001   ;
13'd5113:weight<=16'b0000000000001100   ;
13'd5114:weight<=16'b1111111110110100   ;
13'd5115:weight<=16'b0000000001100001   ;
13'd5116:weight<=16'b0000000010011101   ;
13'd5117:weight<=16'b1111111111110100    ;
13'd5118:weight<=16'b1111111110010011    ;
13'd5119:weight<=16'b0000000000001111    ;
default:weight<=16'd0000000000000000;
endcase
endmodule